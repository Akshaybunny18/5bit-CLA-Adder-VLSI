* SPICE3 file created from Xor.ext - technology: scmos
.include TSMC_180nm.txt
.param LAMBDA = 0.09u
.global gnd vdd
vdd vdd gnd 1.8
.option scale=0.09u

.option scale=0.09u

M1000 gnd a a_156_45# Gnd CMOSN w=40 l=2
+  ad=800 pd=360 as=240 ps=92
M1001 gnd a_94_38# a_236_13# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1002 gnd a_23_6# a_156_n19# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1003 vdd a_94_n26# out w_168_0# CMOSP w=40 l=2
+  ad=960 pd=368 as=400 ps=180
M1004 vdd b a_94_n26# w_88_n32# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1005 a_156_n19# b a_94_n26# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1006 a_23_6# a vdd w_17_0# CMOSP w=40 l=2
+  ad=400 pd=180 as=0 ps=0
M1007 a_236_13# a_94_n26# out Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1008 gnd a a_85_13# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=240 ps=92
M1009 out a_94_38# vdd w_168_0# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 vdd a_23_6# a_94_38# w_88_32# CMOSP w=40 l=2
+  ad=0 pd=0 as=400 ps=180
M1011 a_156_45# a_23_6# a_94_38# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1012 vdd b a_23_6# w_17_0# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1013 a_94_n26# a_23_6# vdd w_88_n32# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
M1014 a_85_13# b a_23_6# Gnd CMOSN w=40 l=2
+  ad=0 pd=0 as=200 ps=90
M1015 a_94_38# a vdd w_88_32# CMOSP w=40 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out gnd 0.07fF
C1 a_94_38# w_88_32# 0.14fF
C2 a_156_45# gnd 0.41fF
C3 b a_94_n26# 0.15fF
C4 vdd w_17_0# 0.06fF
C5 a_94_38# vdd 1.30fF
C6 a w_17_0# 0.08fF
C7 a_94_38# w_168_0# 0.08fF
C8 a_85_13# vdd 0.09fF
C9 a_94_38# a 0.08fF
C10 vdd a_94_n26# 0.90fF
C11 a_156_n19# a_94_n26# 0.45fF
C12 a_94_38# gnd 0.04fF
C13 w_88_n32# a_94_n26# 0.14fF
C14 a_23_6# w_17_0# 0.14fF
C15 a_236_13# gnd 0.41fF
C16 b vdd 0.01fF
C17 w_168_0# a_94_n26# 0.08fF
C18 a_94_38# out 0.08fF
C19 b w_88_n32# 0.08fF
C20 a_85_13# gnd 0.41fF
C21 a_94_38# a_23_6# 0.08fF
C22 a_94_38# a_156_45# 0.41fF
C23 a_236_13# out 0.41fF
C24 gnd a_94_n26# 0.12fF
C25 w_88_32# vdd 0.50fF
C26 b a 0.27fF
C27 a_85_13# a_23_6# 0.41fF
C28 out a_94_n26# 0.08fF
C29 a_23_6# a_94_n26# 0.15fF
C30 w_88_32# a 0.08fF
C31 b a_23_6# 0.40fF
C32 w_88_n32# vdd 0.10fF
C33 w_88_32# a_23_6# 0.08fF
C34 w_168_0# vdd 0.05fF
C35 vdd a 0.33fF
C36 a_156_n19# gnd 0.41fF
C37 vdd gnd 0.10fF
C38 w_88_n32# gnd 0.03fF
C39 vdd out 0.90fF
C40 a_94_38# a_94_n26# 0.31fF
C41 w_168_0# gnd 0.31fF
C42 b w_17_0# 0.08fF
C43 a_23_6# vdd 1.18fF
C44 a_23_6# w_88_n32# 0.08fF
C45 w_168_0# out 0.14fF
C46 a_23_6# a 0.40fF
C47 a_156_n19# Gnd 0.01fF
C48 a_236_13# Gnd 0.01fF
C49 a_94_n26# Gnd 0.45fF
C50 a_85_13# Gnd 0.01fF
C51 b Gnd 0.31fF
C52 a_156_45# Gnd 0.01fF
C53 a_23_6# Gnd 0.43fF
C54 vdd Gnd 0.29fF
C55 gnd Gnd 0.01fF
C56 a Gnd 0.31fF
C57 a_94_38# Gnd 0.41fF
C58 w_88_n32# Gnd 1.67fF
C59 w_168_0# Gnd 1.03fF
C60 w_17_0# Gnd 1.67fF
C61 w_88_32# Gnd 0.02fF

* Testbench for XOR2 gate
* Input signals
Va a gnd 0
Vb b gnd PULSE(0 1.8 15n 0 0 15n 30n)

* Save signals
.save v(a) v(b) v(out)
.tran 50p 160n

.control
run
set curplottitle = "Akshay Chanda 2024102014 - XOR2 Post-Layout"
plot v(b)+3 v(out)

* Propagation delays from b input to output
meas tran tpdr trig v(b) val=0.9 rise=3 targ v(out) val=0.9 rise=3
meas tran tpdf trig v(b) val=0.9 fall=3 targ v(out) val=0.9 fall=3
meas tran tpd param='(tpdr+tpdf)/2'

.endc

.end
