magic
tech scmos
timestamp 1763272488
<< nwell >>
rect 4 36 28 92
<< ntransistor >>
rect 15 8 17 28
<< ptransistor >>
rect 15 42 17 82
<< ndiffusion >>
rect 14 8 15 28
rect 17 8 18 28
<< pdiffusion >>
rect 14 42 15 82
rect 17 42 18 82
<< ndcontact >>
rect 10 8 14 28
rect 18 8 22 28
<< pdcontact >>
rect 10 42 14 82
rect 18 42 22 82
<< polysilicon >>
rect 15 82 17 85
rect 15 28 17 42
rect 15 5 17 8
<< polycontact >>
rect 11 31 15 35
<< metal1 >>
rect 4 88 28 92
rect 10 82 14 88
rect 18 35 22 42
rect 0 31 11 35
rect 18 31 36 35
rect 18 28 22 31
rect 10 4 14 8
rect 4 0 28 4
<< labels >>
rlabel metal1 0 31 4 35 3 in
rlabel metal1 12 0 16 4 1 gnd1
rlabel metal1 32 31 36 35 7 out
rlabel metal1 14 88 18 92 5 vdd1
<< end >>
