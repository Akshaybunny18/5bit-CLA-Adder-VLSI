magic
tech scmos
timestamp 1763233755
<< nwell >>
rect -11 71 21 123
<< ntransistor >>
rect 0 15 2 55
rect 8 15 10 55
<< ptransistor >>
rect 0 77 2 117
rect 8 77 10 117
<< ndiffusion >>
rect -1 15 0 55
rect 2 15 3 55
rect 7 15 8 55
rect 10 15 11 55
<< pdiffusion >>
rect -1 77 0 117
rect 2 77 3 117
rect 7 77 8 117
rect 10 77 11 117
<< ndcontact >>
rect -5 15 -1 55
rect 3 15 7 55
rect 11 15 15 55
<< pdcontact >>
rect -5 77 -1 117
rect 3 77 7 117
rect 11 77 15 117
<< polysilicon >>
rect 0 117 2 130
rect 8 117 10 130
rect 0 55 2 77
rect 8 55 10 77
rect 0 12 2 15
rect 8 12 10 15
<< polycontact >>
rect -1 130 3 134
rect 7 130 11 134
<< metal1 >>
rect -1 134 3 140
rect 7 134 11 140
rect 3 117 7 126
rect -5 73 -1 77
rect 11 73 15 77
rect -5 69 15 73
rect -5 55 -1 69
rect 11 7 15 15
<< labels >>
rlabel metal1 3 122 7 126 1 vdd
rlabel metal1 7 136 11 140 5 b
rlabel metal1 -1 136 3 140 5 a
rlabel metal1 11 7 15 11 1 gnd
rlabel metal1 -5 62 -1 66 1 out
<< end >>
