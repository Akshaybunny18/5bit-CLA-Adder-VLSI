magic
tech scmos
timestamp 1764441304
<< nwell >>
rect -397 79 -364 172
rect -358 93 -334 145
rect -309 93 -283 145
rect -277 79 -253 131
rect -196 78 -163 171
rect -157 92 -133 144
rect -108 92 -82 144
rect -76 78 -52 130
rect 88 64 140 96
rect 383 78 416 171
rect 422 92 446 144
rect 471 92 497 144
rect 503 78 527 130
rect 1127 78 1160 171
rect 1166 92 1190 144
rect 1215 92 1241 144
rect 1247 78 1271 130
rect 17 32 69 64
rect 168 32 220 64
rect 88 0 140 32
rect -396 -114 -363 -21
rect -357 -100 -333 -48
rect -308 -100 -282 -48
rect -276 -114 -252 -62
rect -195 -115 -162 -22
rect 88 -38 140 -6
rect -156 -101 -132 -49
rect -107 -101 -81 -49
rect -75 -115 -51 -63
rect 88 -85 140 -53
rect 215 -55 267 -31
rect 390 -62 442 -30
rect 845 -36 897 -4
rect 557 -70 609 -38
rect 774 -68 826 -36
rect 925 -68 977 -36
rect 17 -117 69 -85
rect 168 -117 220 -85
rect 845 -100 897 -68
rect 88 -149 140 -117
rect 88 -187 140 -155
rect 391 -165 443 -125
rect -398 -302 -365 -209
rect -359 -288 -335 -236
rect -310 -288 -284 -236
rect -278 -302 -254 -250
rect -197 -303 -164 -210
rect 88 -235 140 -203
rect 215 -204 267 -180
rect 390 -206 442 -174
rect 580 -181 632 -141
rect 845 -145 897 -113
rect 1128 -115 1161 -22
rect 1167 -101 1191 -49
rect 1216 -101 1242 -49
rect 1248 -115 1272 -63
rect 774 -177 826 -145
rect 925 -177 977 -145
rect 845 -209 897 -177
rect -158 -289 -134 -237
rect -109 -289 -83 -237
rect -77 -303 -53 -251
rect 17 -267 69 -235
rect 168 -267 220 -235
rect 88 -299 140 -267
rect 390 -290 442 -242
rect 845 -255 897 -223
rect 774 -287 826 -255
rect 925 -287 977 -255
rect 88 -337 140 -305
rect 88 -384 140 -352
rect 214 -354 266 -330
rect 391 -336 443 -296
rect 390 -377 442 -345
rect 570 -351 622 -303
rect 845 -319 897 -287
rect 1126 -303 1159 -210
rect 1165 -289 1189 -237
rect 1214 -289 1240 -237
rect 1246 -303 1270 -251
rect 845 -366 897 -334
rect -397 -493 -364 -400
rect -358 -479 -334 -427
rect -309 -479 -283 -427
rect -277 -493 -253 -441
rect -196 -494 -163 -401
rect 17 -416 69 -384
rect 168 -416 220 -384
rect 774 -398 826 -366
rect 925 -398 977 -366
rect -157 -480 -133 -428
rect -108 -480 -82 -428
rect -76 -494 -52 -442
rect 88 -448 140 -416
rect 88 -486 140 -454
rect 390 -472 442 -416
rect 845 -430 897 -398
rect 88 -534 140 -502
rect 214 -503 266 -479
rect 390 -527 442 -479
rect 1127 -494 1160 -401
rect 1166 -480 1190 -428
rect 1215 -480 1241 -428
rect 1247 -494 1271 -442
rect 17 -566 69 -534
rect 168 -566 220 -534
rect -395 -683 -362 -590
rect -356 -669 -332 -617
rect -307 -669 -281 -617
rect -275 -683 -251 -631
rect -194 -684 -161 -591
rect 88 -598 140 -566
rect 391 -573 443 -533
rect -155 -670 -131 -618
rect -106 -670 -80 -618
rect -74 -684 -50 -632
rect 88 -636 140 -604
rect 390 -614 442 -582
rect 546 -607 598 -551
rect 214 -653 266 -629
rect 1129 -684 1162 -591
rect 1168 -670 1192 -618
rect 1217 -670 1243 -618
rect 1249 -684 1273 -632
<< ntransistor >>
rect -386 30 -384 50
rect -347 44 -345 84
rect -339 44 -337 84
rect -298 44 -296 84
rect -290 44 -288 84
rect -266 51 -264 71
rect -185 29 -183 49
rect -146 43 -144 83
rect -138 43 -136 83
rect -97 43 -95 83
rect -89 43 -87 83
rect 156 83 196 85
rect 156 75 196 77
rect -65 50 -63 70
rect 85 51 125 53
rect 236 51 276 53
rect 85 43 125 45
rect 236 43 276 45
rect 394 29 396 49
rect 433 43 435 83
rect 441 43 443 83
rect 482 43 484 83
rect 490 43 492 83
rect 514 50 516 70
rect 1138 29 1140 49
rect 1177 43 1179 83
rect 1185 43 1187 83
rect 1226 43 1228 83
rect 1234 43 1236 83
rect 1258 50 1260 70
rect 156 19 196 21
rect 156 11 196 13
rect 156 -19 196 -17
rect 913 -17 953 -15
rect 156 -27 196 -25
rect 913 -25 953 -23
rect 275 -44 295 -42
rect 458 -43 498 -41
rect 458 -51 498 -49
rect 625 -51 665 -49
rect 842 -49 882 -47
rect 625 -59 665 -57
rect 993 -49 1033 -47
rect 842 -57 882 -55
rect 993 -57 1033 -55
rect 156 -66 196 -64
rect -385 -163 -383 -143
rect -346 -149 -344 -109
rect -338 -149 -336 -109
rect -297 -149 -295 -109
rect -289 -149 -287 -109
rect 156 -74 196 -72
rect 913 -81 953 -79
rect 913 -89 953 -87
rect 85 -98 125 -96
rect 236 -98 276 -96
rect 85 -106 125 -104
rect -265 -142 -263 -122
rect -184 -164 -182 -144
rect -145 -150 -143 -110
rect -137 -150 -135 -110
rect -96 -150 -94 -110
rect -88 -150 -86 -110
rect 236 -106 276 -104
rect -64 -143 -62 -123
rect 913 -126 953 -124
rect 156 -130 196 -128
rect 156 -138 196 -136
rect 913 -134 953 -132
rect 453 -138 513 -136
rect 453 -146 513 -144
rect 453 -154 513 -152
rect 642 -154 702 -152
rect 842 -158 882 -156
rect 642 -162 702 -160
rect 156 -168 196 -166
rect 993 -158 1033 -156
rect 842 -166 882 -164
rect 642 -170 702 -168
rect 156 -176 196 -174
rect 1139 -164 1141 -144
rect 1178 -150 1180 -110
rect 1186 -150 1188 -110
rect 1227 -150 1229 -110
rect 1235 -150 1237 -110
rect 1259 -143 1261 -123
rect 993 -166 1033 -164
rect 458 -187 498 -185
rect 275 -193 295 -191
rect 913 -190 953 -188
rect 458 -195 498 -193
rect 913 -198 953 -196
rect 156 -216 196 -214
rect 156 -224 196 -222
rect 913 -236 953 -234
rect 85 -248 125 -246
rect 913 -244 953 -242
rect 236 -248 276 -246
rect 85 -256 125 -254
rect -387 -351 -385 -331
rect -348 -337 -346 -297
rect -340 -337 -338 -297
rect -299 -337 -297 -297
rect -291 -337 -289 -297
rect 236 -256 276 -254
rect 452 -255 532 -253
rect 452 -263 532 -261
rect 842 -268 882 -266
rect 452 -271 532 -269
rect 156 -280 196 -278
rect 993 -268 1033 -266
rect 842 -276 882 -274
rect 452 -279 532 -277
rect 993 -276 1033 -274
rect 156 -288 196 -286
rect -267 -330 -265 -310
rect -186 -352 -184 -332
rect -147 -338 -145 -298
rect -139 -338 -137 -298
rect -98 -338 -96 -298
rect -90 -338 -88 -298
rect 913 -300 953 -298
rect 453 -309 513 -307
rect 913 -308 953 -306
rect -66 -331 -64 -311
rect 156 -318 196 -316
rect 453 -317 513 -315
rect 632 -316 712 -314
rect 156 -326 196 -324
rect 453 -325 513 -323
rect 632 -324 712 -322
rect 632 -332 712 -330
rect 632 -340 712 -338
rect 274 -343 294 -341
rect 913 -347 953 -345
rect 1137 -352 1139 -332
rect 1176 -338 1178 -298
rect 1184 -338 1186 -298
rect 1225 -338 1227 -298
rect 1233 -338 1235 -298
rect 1257 -331 1259 -311
rect 913 -355 953 -353
rect 458 -358 498 -356
rect 156 -365 196 -363
rect 458 -366 498 -364
rect 156 -373 196 -371
rect 842 -379 882 -377
rect 993 -379 1033 -377
rect 842 -387 882 -385
rect 85 -397 125 -395
rect 993 -387 1033 -385
rect 236 -397 276 -395
rect 85 -405 125 -403
rect 236 -405 276 -403
rect 913 -411 953 -409
rect 913 -419 953 -417
rect 156 -429 196 -427
rect 452 -429 552 -427
rect 156 -437 196 -435
rect 452 -437 552 -435
rect 452 -445 552 -443
rect -386 -542 -384 -522
rect -347 -528 -345 -488
rect -339 -528 -337 -488
rect -298 -528 -296 -488
rect -290 -528 -288 -488
rect 452 -453 552 -451
rect 452 -461 552 -459
rect 156 -467 196 -465
rect 156 -475 196 -473
rect -266 -521 -264 -501
rect -185 -543 -183 -523
rect -146 -529 -144 -489
rect -138 -529 -136 -489
rect -97 -529 -95 -489
rect -89 -529 -87 -489
rect 274 -492 294 -490
rect 452 -492 532 -490
rect 452 -500 532 -498
rect -65 -522 -63 -502
rect 452 -508 532 -506
rect 156 -515 196 -513
rect 452 -516 532 -514
rect 156 -523 196 -521
rect 85 -547 125 -545
rect 236 -547 276 -545
rect 1138 -543 1140 -523
rect 1177 -529 1179 -489
rect 1185 -529 1187 -489
rect 1226 -529 1228 -489
rect 1234 -529 1236 -489
rect 1258 -522 1260 -502
rect 453 -546 513 -544
rect 85 -555 125 -553
rect 236 -555 276 -553
rect 453 -554 513 -552
rect 453 -562 513 -560
rect 608 -564 708 -562
rect 608 -572 708 -570
rect 156 -579 196 -577
rect 608 -580 708 -578
rect 156 -587 196 -585
rect 608 -588 708 -586
rect 458 -595 498 -593
rect 608 -596 708 -594
rect 458 -603 498 -601
rect 156 -617 196 -615
rect 156 -625 196 -623
rect -384 -732 -382 -712
rect -345 -718 -343 -678
rect -337 -718 -335 -678
rect -296 -718 -294 -678
rect -288 -718 -286 -678
rect 274 -642 294 -640
rect -264 -711 -262 -691
rect -183 -733 -181 -713
rect -144 -719 -142 -679
rect -136 -719 -134 -679
rect -95 -719 -93 -679
rect -87 -719 -85 -679
rect -63 -712 -61 -692
rect 1140 -733 1142 -713
rect 1179 -719 1181 -679
rect 1187 -719 1189 -679
rect 1228 -719 1230 -679
rect 1236 -719 1238 -679
rect 1260 -712 1262 -692
<< ptransistor >>
rect -386 86 -384 166
rect -378 86 -376 166
rect -347 99 -345 139
rect -298 99 -296 139
rect -266 85 -264 125
rect -185 85 -183 165
rect -177 85 -175 165
rect -146 98 -144 138
rect -97 98 -95 138
rect -65 84 -63 124
rect 394 85 396 165
rect 402 85 404 165
rect 433 98 435 138
rect 482 98 484 138
rect 94 83 134 85
rect 94 75 134 77
rect 514 84 516 124
rect 1138 85 1140 165
rect 1146 85 1148 165
rect 1177 98 1179 138
rect 1226 98 1228 138
rect 23 51 63 53
rect 174 51 214 53
rect 23 43 63 45
rect 174 43 214 45
rect 1258 84 1260 124
rect 94 19 134 21
rect 94 11 134 13
rect -385 -107 -383 -27
rect -377 -107 -375 -27
rect 94 -19 134 -17
rect 851 -17 891 -15
rect 94 -27 134 -25
rect 851 -25 891 -23
rect -346 -94 -344 -54
rect -297 -94 -295 -54
rect -265 -108 -263 -68
rect -184 -108 -182 -28
rect -176 -108 -174 -28
rect 221 -44 261 -42
rect 396 -43 436 -41
rect 396 -51 436 -49
rect -145 -95 -143 -55
rect -96 -95 -94 -55
rect 563 -51 603 -49
rect 780 -49 820 -47
rect 563 -59 603 -57
rect 931 -49 971 -47
rect 780 -57 820 -55
rect 931 -57 971 -55
rect 94 -66 134 -64
rect -64 -109 -62 -69
rect 94 -74 134 -72
rect 851 -81 891 -79
rect 851 -89 891 -87
rect 23 -98 63 -96
rect 174 -98 214 -96
rect 23 -106 63 -104
rect 174 -106 214 -104
rect 1139 -108 1141 -28
rect 1147 -108 1149 -28
rect 1178 -95 1180 -55
rect 1227 -95 1229 -55
rect 1259 -109 1261 -69
rect 851 -126 891 -124
rect 94 -130 134 -128
rect 94 -138 134 -136
rect 851 -134 891 -132
rect 397 -138 437 -136
rect 397 -146 437 -144
rect 397 -154 437 -152
rect 586 -154 626 -152
rect 780 -158 820 -156
rect 586 -162 626 -160
rect 94 -168 134 -166
rect 931 -158 971 -156
rect 780 -166 820 -164
rect 586 -170 626 -168
rect 94 -176 134 -174
rect 931 -166 971 -164
rect 396 -187 436 -185
rect 221 -193 261 -191
rect 851 -190 891 -188
rect 396 -195 436 -193
rect 851 -198 891 -196
rect -387 -295 -385 -215
rect -379 -295 -377 -215
rect -348 -282 -346 -242
rect -299 -282 -297 -242
rect -267 -296 -265 -256
rect -186 -296 -184 -216
rect -178 -296 -176 -216
rect 94 -216 134 -214
rect 94 -224 134 -222
rect 851 -236 891 -234
rect -147 -283 -145 -243
rect -98 -283 -96 -243
rect 23 -248 63 -246
rect 851 -244 891 -242
rect 174 -248 214 -246
rect 23 -256 63 -254
rect -66 -297 -64 -257
rect 174 -256 214 -254
rect 396 -255 436 -253
rect 396 -263 436 -261
rect 780 -268 820 -266
rect 396 -271 436 -269
rect 94 -280 134 -278
rect 931 -268 971 -266
rect 780 -276 820 -274
rect 396 -279 436 -277
rect 931 -276 971 -274
rect 94 -288 134 -286
rect 1137 -296 1139 -216
rect 1145 -296 1147 -216
rect 1176 -283 1178 -243
rect 1225 -283 1227 -243
rect 851 -300 891 -298
rect 397 -309 437 -307
rect 851 -308 891 -306
rect 1257 -297 1259 -257
rect 94 -318 134 -316
rect 397 -317 437 -315
rect 576 -316 616 -314
rect 94 -326 134 -324
rect 397 -325 437 -323
rect 576 -324 616 -322
rect 576 -332 616 -330
rect 576 -340 616 -338
rect 220 -343 260 -341
rect 851 -347 891 -345
rect 851 -355 891 -353
rect 396 -358 436 -356
rect 94 -365 134 -363
rect 396 -366 436 -364
rect 94 -373 134 -371
rect 780 -379 820 -377
rect 931 -379 971 -377
rect 780 -387 820 -385
rect -386 -486 -384 -406
rect -378 -486 -376 -406
rect 23 -397 63 -395
rect 931 -387 971 -385
rect 174 -397 214 -395
rect 23 -405 63 -403
rect -347 -473 -345 -433
rect -298 -473 -296 -433
rect -266 -487 -264 -447
rect -185 -487 -183 -407
rect -177 -487 -175 -407
rect 174 -405 214 -403
rect 851 -411 891 -409
rect 851 -419 891 -417
rect 94 -429 134 -427
rect -146 -474 -144 -434
rect -97 -474 -95 -434
rect 396 -429 436 -427
rect 94 -437 134 -435
rect 396 -437 436 -435
rect 396 -445 436 -443
rect -65 -488 -63 -448
rect 396 -453 436 -451
rect 396 -461 436 -459
rect 94 -467 134 -465
rect 94 -475 134 -473
rect 220 -492 260 -490
rect 1138 -487 1140 -407
rect 1146 -487 1148 -407
rect 1177 -474 1179 -434
rect 1226 -474 1228 -434
rect 396 -492 436 -490
rect 396 -500 436 -498
rect 1258 -488 1260 -448
rect 396 -508 436 -506
rect 94 -515 134 -513
rect 396 -516 436 -514
rect 94 -523 134 -521
rect 23 -547 63 -545
rect 174 -547 214 -545
rect 397 -546 437 -544
rect 23 -555 63 -553
rect 174 -555 214 -553
rect 397 -554 437 -552
rect 397 -562 437 -560
rect 552 -564 592 -562
rect 552 -572 592 -570
rect 94 -579 134 -577
rect -384 -676 -382 -596
rect -376 -676 -374 -596
rect 552 -580 592 -578
rect 94 -587 134 -585
rect 552 -588 592 -586
rect 396 -595 436 -593
rect -345 -663 -343 -623
rect -296 -663 -294 -623
rect -264 -677 -262 -637
rect -183 -677 -181 -597
rect -175 -677 -173 -597
rect 552 -596 592 -594
rect 396 -603 436 -601
rect 94 -617 134 -615
rect -144 -664 -142 -624
rect -95 -664 -93 -624
rect 94 -625 134 -623
rect -63 -678 -61 -638
rect 220 -642 260 -640
rect 1140 -677 1142 -597
rect 1148 -677 1150 -597
rect 1179 -664 1181 -624
rect 1228 -664 1230 -624
rect 1260 -678 1262 -638
<< ndiffusion >>
rect -387 30 -386 50
rect -384 30 -383 50
rect -348 44 -347 84
rect -345 44 -344 84
rect -340 44 -339 84
rect -337 44 -336 84
rect -299 44 -298 84
rect -296 44 -295 84
rect -291 44 -290 84
rect -288 44 -287 84
rect -267 51 -266 71
rect -264 51 -263 71
rect -186 29 -185 49
rect -183 29 -182 49
rect -147 43 -146 83
rect -144 43 -143 83
rect -139 43 -138 83
rect -136 43 -135 83
rect -98 43 -97 83
rect -95 43 -94 83
rect -90 43 -89 83
rect -87 43 -86 83
rect 156 85 196 86
rect 156 82 196 83
rect 156 77 196 78
rect 156 74 196 75
rect -66 50 -65 70
rect -63 50 -62 70
rect 85 53 125 54
rect 85 50 125 51
rect 236 53 276 54
rect 85 45 125 46
rect 85 42 125 43
rect 236 50 276 51
rect 236 45 276 46
rect 236 42 276 43
rect 393 29 394 49
rect 396 29 397 49
rect 432 43 433 83
rect 435 43 436 83
rect 440 43 441 83
rect 443 43 444 83
rect 481 43 482 83
rect 484 43 485 83
rect 489 43 490 83
rect 492 43 493 83
rect 513 50 514 70
rect 516 50 517 70
rect 1137 29 1138 49
rect 1140 29 1141 49
rect 1176 43 1177 83
rect 1179 43 1180 83
rect 1184 43 1185 83
rect 1187 43 1188 83
rect 1225 43 1226 83
rect 1228 43 1229 83
rect 1233 43 1234 83
rect 1236 43 1237 83
rect 1257 50 1258 70
rect 1260 50 1261 70
rect 156 21 196 22
rect 156 18 196 19
rect 156 13 196 14
rect 156 10 196 11
rect 156 -17 196 -16
rect 913 -15 953 -14
rect 156 -20 196 -19
rect 156 -25 196 -24
rect 913 -18 953 -17
rect 913 -23 953 -22
rect 156 -28 196 -27
rect 913 -26 953 -25
rect 275 -42 295 -41
rect 458 -41 498 -40
rect 275 -45 295 -44
rect 458 -44 498 -43
rect 458 -49 498 -48
rect 458 -52 498 -51
rect 625 -49 665 -48
rect 842 -47 882 -46
rect 625 -52 665 -51
rect 625 -57 665 -56
rect 842 -50 882 -49
rect 993 -47 1033 -46
rect 842 -55 882 -54
rect 156 -64 196 -63
rect 625 -60 665 -59
rect 842 -58 882 -57
rect 993 -50 1033 -49
rect 993 -55 1033 -54
rect 993 -58 1033 -57
rect -386 -163 -385 -143
rect -383 -163 -382 -143
rect -347 -149 -346 -109
rect -344 -149 -343 -109
rect -339 -149 -338 -109
rect -336 -149 -335 -109
rect -298 -149 -297 -109
rect -295 -149 -294 -109
rect -290 -149 -289 -109
rect -287 -149 -286 -109
rect 156 -67 196 -66
rect 156 -72 196 -71
rect 156 -75 196 -74
rect 913 -79 953 -78
rect 913 -82 953 -81
rect 913 -87 953 -86
rect 85 -96 125 -95
rect 85 -99 125 -98
rect 913 -90 953 -89
rect 236 -96 276 -95
rect 85 -104 125 -103
rect -266 -142 -265 -122
rect -263 -142 -262 -122
rect -185 -164 -184 -144
rect -182 -164 -181 -144
rect -146 -150 -145 -110
rect -143 -150 -142 -110
rect -138 -150 -137 -110
rect -135 -150 -134 -110
rect -97 -150 -96 -110
rect -94 -150 -93 -110
rect -89 -150 -88 -110
rect -86 -150 -85 -110
rect 85 -107 125 -106
rect 236 -99 276 -98
rect 236 -104 276 -103
rect 236 -107 276 -106
rect -65 -143 -64 -123
rect -62 -143 -61 -123
rect 913 -124 953 -123
rect 156 -128 196 -127
rect 156 -131 196 -130
rect 156 -136 196 -135
rect 156 -139 196 -138
rect 913 -127 953 -126
rect 913 -132 953 -131
rect 453 -136 513 -135
rect 453 -139 513 -138
rect 913 -135 953 -134
rect 453 -144 513 -143
rect 453 -147 513 -146
rect 453 -152 513 -151
rect 453 -155 513 -154
rect 642 -152 702 -151
rect 642 -155 702 -154
rect 842 -156 882 -155
rect 642 -160 702 -159
rect 156 -166 196 -165
rect 156 -169 196 -168
rect 642 -163 702 -162
rect 842 -159 882 -158
rect 993 -156 1033 -155
rect 842 -164 882 -163
rect 642 -168 702 -167
rect 156 -174 196 -173
rect 642 -171 702 -170
rect 842 -167 882 -166
rect 993 -159 1033 -158
rect 993 -164 1033 -163
rect 1138 -164 1139 -144
rect 1141 -164 1142 -144
rect 1177 -150 1178 -110
rect 1180 -150 1181 -110
rect 1185 -150 1186 -110
rect 1188 -150 1189 -110
rect 1226 -150 1227 -110
rect 1229 -150 1230 -110
rect 1234 -150 1235 -110
rect 1237 -150 1238 -110
rect 1258 -143 1259 -123
rect 1261 -143 1262 -123
rect 993 -167 1033 -166
rect 156 -177 196 -176
rect 458 -185 498 -184
rect 275 -191 295 -190
rect 275 -194 295 -193
rect 458 -188 498 -187
rect 913 -188 953 -187
rect 458 -193 498 -192
rect 458 -196 498 -195
rect 913 -191 953 -190
rect 913 -196 953 -195
rect 913 -199 953 -198
rect 156 -214 196 -213
rect 156 -217 196 -216
rect 156 -222 196 -221
rect 156 -225 196 -224
rect 913 -234 953 -233
rect 85 -246 125 -245
rect 85 -249 125 -248
rect 913 -237 953 -236
rect 913 -242 953 -241
rect 236 -246 276 -245
rect 85 -254 125 -253
rect -388 -351 -387 -331
rect -385 -351 -384 -331
rect -349 -337 -348 -297
rect -346 -337 -345 -297
rect -341 -337 -340 -297
rect -338 -337 -337 -297
rect -300 -337 -299 -297
rect -297 -337 -296 -297
rect -292 -337 -291 -297
rect -289 -337 -288 -297
rect 85 -257 125 -256
rect 236 -249 276 -248
rect 236 -254 276 -253
rect 913 -245 953 -244
rect 452 -253 532 -252
rect 236 -257 276 -256
rect 452 -256 532 -255
rect 452 -261 532 -260
rect 452 -264 532 -263
rect 452 -269 532 -268
rect 842 -266 882 -265
rect 156 -278 196 -277
rect 452 -272 532 -271
rect 452 -277 532 -276
rect 842 -269 882 -268
rect 993 -266 1033 -265
rect 842 -274 882 -273
rect 156 -281 196 -280
rect 452 -280 532 -279
rect 842 -277 882 -276
rect 993 -269 1033 -268
rect 993 -274 1033 -273
rect 993 -277 1033 -276
rect 156 -286 196 -285
rect 156 -289 196 -288
rect -268 -330 -267 -310
rect -265 -330 -264 -310
rect -187 -352 -186 -332
rect -184 -352 -183 -332
rect -148 -338 -147 -298
rect -145 -338 -144 -298
rect -140 -338 -139 -298
rect -137 -338 -136 -298
rect -99 -338 -98 -298
rect -96 -338 -95 -298
rect -91 -338 -90 -298
rect -88 -338 -87 -298
rect 913 -298 953 -297
rect 453 -307 513 -306
rect 913 -301 953 -300
rect 913 -306 953 -305
rect -67 -331 -66 -311
rect -64 -331 -63 -311
rect 156 -316 196 -315
rect 453 -310 513 -309
rect 453 -315 513 -314
rect 913 -309 953 -308
rect 632 -314 712 -313
rect 156 -319 196 -318
rect 156 -324 196 -323
rect 453 -318 513 -317
rect 453 -323 513 -322
rect 632 -317 712 -316
rect 632 -322 712 -321
rect 156 -327 196 -326
rect 453 -326 513 -325
rect 632 -325 712 -324
rect 632 -330 712 -329
rect 274 -341 294 -340
rect 632 -333 712 -332
rect 632 -338 712 -337
rect 274 -344 294 -343
rect 632 -341 712 -340
rect 913 -345 953 -344
rect 458 -356 498 -355
rect 913 -348 953 -347
rect 1136 -352 1137 -332
rect 1139 -352 1140 -332
rect 1175 -338 1176 -298
rect 1178 -338 1179 -298
rect 1183 -338 1184 -298
rect 1186 -338 1187 -298
rect 1224 -338 1225 -298
rect 1227 -338 1228 -298
rect 1232 -338 1233 -298
rect 1235 -338 1236 -298
rect 1256 -331 1257 -311
rect 1259 -331 1260 -311
rect 913 -353 953 -352
rect 156 -363 196 -362
rect 156 -366 196 -365
rect 458 -359 498 -358
rect 913 -356 953 -355
rect 458 -364 498 -363
rect 156 -371 196 -370
rect 458 -367 498 -366
rect 156 -374 196 -373
rect 842 -377 882 -376
rect 842 -380 882 -379
rect 993 -377 1033 -376
rect 842 -385 882 -384
rect 85 -395 125 -394
rect 85 -398 125 -397
rect 842 -388 882 -387
rect 993 -380 1033 -379
rect 993 -385 1033 -384
rect 993 -388 1033 -387
rect 236 -395 276 -394
rect 85 -403 125 -402
rect 85 -406 125 -405
rect 236 -398 276 -397
rect 236 -403 276 -402
rect 236 -406 276 -405
rect 913 -409 953 -408
rect 913 -412 953 -411
rect 913 -417 953 -416
rect 156 -427 196 -426
rect 156 -430 196 -429
rect 913 -420 953 -419
rect 452 -427 552 -426
rect 156 -435 196 -434
rect 156 -438 196 -437
rect 452 -430 552 -429
rect 452 -435 552 -434
rect 452 -438 552 -437
rect 452 -443 552 -442
rect -387 -542 -386 -522
rect -384 -542 -383 -522
rect -348 -528 -347 -488
rect -345 -528 -344 -488
rect -340 -528 -339 -488
rect -337 -528 -336 -488
rect -299 -528 -298 -488
rect -296 -528 -295 -488
rect -291 -528 -290 -488
rect -288 -528 -287 -488
rect 452 -446 552 -445
rect 452 -451 552 -450
rect 452 -454 552 -453
rect 452 -459 552 -458
rect 156 -465 196 -464
rect 452 -462 552 -461
rect 156 -468 196 -467
rect 156 -473 196 -472
rect 156 -476 196 -475
rect -267 -521 -266 -501
rect -264 -521 -263 -501
rect -186 -543 -185 -523
rect -183 -543 -182 -523
rect -147 -529 -146 -489
rect -144 -529 -143 -489
rect -139 -529 -138 -489
rect -136 -529 -135 -489
rect -98 -529 -97 -489
rect -95 -529 -94 -489
rect -90 -529 -89 -489
rect -87 -529 -86 -489
rect 274 -490 294 -489
rect 274 -493 294 -492
rect 452 -490 532 -489
rect 452 -493 532 -492
rect 452 -498 532 -497
rect -66 -522 -65 -502
rect -63 -522 -62 -502
rect 452 -501 532 -500
rect 452 -506 532 -505
rect 156 -513 196 -512
rect 156 -516 196 -515
rect 452 -509 532 -508
rect 452 -514 532 -513
rect 156 -521 196 -520
rect 452 -517 532 -516
rect 156 -524 196 -523
rect 85 -545 125 -544
rect 85 -548 125 -547
rect 236 -545 276 -544
rect 1137 -543 1138 -523
rect 1140 -543 1141 -523
rect 1176 -529 1177 -489
rect 1179 -529 1180 -489
rect 1184 -529 1185 -489
rect 1187 -529 1188 -489
rect 1225 -529 1226 -489
rect 1228 -529 1229 -489
rect 1233 -529 1234 -489
rect 1236 -529 1237 -489
rect 1257 -522 1258 -502
rect 1260 -522 1261 -502
rect 453 -544 513 -543
rect 85 -553 125 -552
rect 85 -556 125 -555
rect 236 -548 276 -547
rect 236 -553 276 -552
rect 453 -547 513 -546
rect 453 -552 513 -551
rect 236 -556 276 -555
rect 453 -555 513 -554
rect 453 -560 513 -559
rect 453 -563 513 -562
rect 608 -562 708 -561
rect 608 -565 708 -564
rect 608 -570 708 -569
rect 156 -577 196 -576
rect 156 -580 196 -579
rect 608 -573 708 -572
rect 608 -578 708 -577
rect 156 -585 196 -584
rect 156 -588 196 -587
rect 608 -581 708 -580
rect 608 -586 708 -585
rect 458 -593 498 -592
rect 458 -596 498 -595
rect 608 -589 708 -588
rect 608 -594 708 -593
rect 458 -601 498 -600
rect 608 -597 708 -596
rect 458 -604 498 -603
rect 156 -615 196 -614
rect 156 -618 196 -617
rect 156 -623 196 -622
rect 156 -626 196 -625
rect -385 -732 -384 -712
rect -382 -732 -381 -712
rect -346 -718 -345 -678
rect -343 -718 -342 -678
rect -338 -718 -337 -678
rect -335 -718 -334 -678
rect -297 -718 -296 -678
rect -294 -718 -293 -678
rect -289 -718 -288 -678
rect -286 -718 -285 -678
rect 274 -640 294 -639
rect 274 -643 294 -642
rect -265 -711 -264 -691
rect -262 -711 -261 -691
rect -184 -733 -183 -713
rect -181 -733 -180 -713
rect -145 -719 -144 -679
rect -142 -719 -141 -679
rect -137 -719 -136 -679
rect -134 -719 -133 -679
rect -96 -719 -95 -679
rect -93 -719 -92 -679
rect -88 -719 -87 -679
rect -85 -719 -84 -679
rect -64 -712 -63 -692
rect -61 -712 -60 -692
rect 1139 -733 1140 -713
rect 1142 -733 1143 -713
rect 1178 -719 1179 -679
rect 1181 -719 1182 -679
rect 1186 -719 1187 -679
rect 1189 -719 1190 -679
rect 1227 -719 1228 -679
rect 1230 -719 1231 -679
rect 1235 -719 1236 -679
rect 1238 -719 1239 -679
rect 1259 -712 1260 -692
rect 1262 -712 1263 -692
<< pdiffusion >>
rect -387 86 -386 166
rect -384 86 -383 166
rect -379 86 -378 166
rect -376 86 -375 166
rect -371 86 -370 166
rect -348 99 -347 139
rect -345 99 -344 139
rect -299 99 -298 139
rect -296 99 -295 139
rect -267 85 -266 125
rect -264 85 -263 125
rect -186 85 -185 165
rect -183 85 -182 165
rect -178 85 -177 165
rect -175 85 -174 165
rect -170 85 -169 165
rect -147 98 -146 138
rect -144 98 -143 138
rect -98 98 -97 138
rect -95 98 -94 138
rect -66 84 -65 124
rect -63 84 -62 124
rect 94 85 134 86
rect 393 85 394 165
rect 396 85 397 165
rect 401 85 402 165
rect 404 85 405 165
rect 409 85 410 165
rect 432 98 433 138
rect 435 98 436 138
rect 481 98 482 138
rect 484 98 485 138
rect 94 82 134 83
rect 94 77 134 78
rect 94 74 134 75
rect 513 84 514 124
rect 516 84 517 124
rect 1137 85 1138 165
rect 1140 85 1141 165
rect 1145 85 1146 165
rect 1148 85 1149 165
rect 1153 85 1154 165
rect 1176 98 1177 138
rect 1179 98 1180 138
rect 1225 98 1226 138
rect 1228 98 1229 138
rect 23 53 63 54
rect 23 50 63 51
rect 23 45 63 46
rect 174 53 214 54
rect 174 50 214 51
rect 23 42 63 43
rect 174 45 214 46
rect 174 42 214 43
rect 1257 84 1258 124
rect 1260 84 1261 124
rect 94 21 134 22
rect 94 18 134 19
rect 94 13 134 14
rect 94 10 134 11
rect -386 -107 -385 -27
rect -383 -107 -382 -27
rect -378 -107 -377 -27
rect -375 -107 -374 -27
rect -370 -107 -369 -27
rect 94 -17 134 -16
rect 851 -15 891 -14
rect 851 -18 891 -17
rect 94 -20 134 -19
rect 94 -25 134 -24
rect 851 -23 891 -22
rect 851 -26 891 -25
rect 94 -28 134 -27
rect -347 -94 -346 -54
rect -344 -94 -343 -54
rect -298 -94 -297 -54
rect -295 -94 -294 -54
rect -266 -108 -265 -68
rect -263 -108 -262 -68
rect -185 -108 -184 -28
rect -182 -108 -181 -28
rect -177 -108 -176 -28
rect -174 -108 -173 -28
rect -169 -108 -168 -28
rect 221 -42 261 -41
rect 396 -41 436 -40
rect 396 -44 436 -43
rect 221 -45 261 -44
rect 396 -49 436 -48
rect 396 -52 436 -51
rect -146 -95 -145 -55
rect -143 -95 -142 -55
rect -97 -95 -96 -55
rect -94 -95 -93 -55
rect 563 -49 603 -48
rect 780 -47 820 -46
rect 780 -50 820 -49
rect 563 -52 603 -51
rect 94 -64 134 -63
rect 563 -57 603 -56
rect 780 -55 820 -54
rect 931 -47 971 -46
rect 931 -50 971 -49
rect 780 -58 820 -57
rect 563 -60 603 -59
rect 931 -55 971 -54
rect 931 -58 971 -57
rect 94 -67 134 -66
rect -65 -109 -64 -69
rect -62 -109 -61 -69
rect 94 -72 134 -71
rect 94 -75 134 -74
rect 851 -79 891 -78
rect 851 -82 891 -81
rect 851 -87 891 -86
rect 851 -90 891 -89
rect 23 -96 63 -95
rect 23 -99 63 -98
rect 23 -104 63 -103
rect 174 -96 214 -95
rect 174 -99 214 -98
rect 23 -107 63 -106
rect 174 -104 214 -103
rect 174 -107 214 -106
rect 1138 -108 1139 -28
rect 1141 -108 1142 -28
rect 1146 -108 1147 -28
rect 1149 -108 1150 -28
rect 1154 -108 1155 -28
rect 1177 -95 1178 -55
rect 1180 -95 1181 -55
rect 1226 -95 1227 -55
rect 1229 -95 1230 -55
rect 1258 -109 1259 -69
rect 1261 -109 1262 -69
rect 94 -128 134 -127
rect 851 -124 891 -123
rect 851 -127 891 -126
rect 94 -131 134 -130
rect 94 -136 134 -135
rect 94 -139 134 -138
rect 397 -136 437 -135
rect 851 -132 891 -131
rect 851 -135 891 -134
rect 397 -139 437 -138
rect 397 -144 437 -143
rect 397 -147 437 -146
rect 397 -152 437 -151
rect 397 -155 437 -154
rect 586 -152 626 -151
rect 586 -155 626 -154
rect 94 -166 134 -165
rect 586 -160 626 -159
rect 780 -156 820 -155
rect 780 -159 820 -158
rect 586 -163 626 -162
rect 94 -169 134 -168
rect 94 -174 134 -173
rect 586 -168 626 -167
rect 780 -164 820 -163
rect 931 -156 971 -155
rect 931 -159 971 -158
rect 780 -167 820 -166
rect 586 -171 626 -170
rect 931 -164 971 -163
rect 931 -167 971 -166
rect 94 -177 134 -176
rect 221 -191 261 -190
rect 396 -185 436 -184
rect 396 -188 436 -187
rect 221 -194 261 -193
rect 396 -193 436 -192
rect 851 -188 891 -187
rect 851 -191 891 -190
rect 396 -196 436 -195
rect 851 -196 891 -195
rect 851 -199 891 -198
rect -388 -295 -387 -215
rect -385 -295 -384 -215
rect -380 -295 -379 -215
rect -377 -295 -376 -215
rect -372 -295 -371 -215
rect -349 -282 -348 -242
rect -346 -282 -345 -242
rect -300 -282 -299 -242
rect -297 -282 -296 -242
rect -268 -296 -267 -256
rect -265 -296 -264 -256
rect -187 -296 -186 -216
rect -184 -296 -183 -216
rect -179 -296 -178 -216
rect -176 -296 -175 -216
rect -171 -296 -170 -216
rect 94 -214 134 -213
rect 94 -217 134 -216
rect 94 -222 134 -221
rect 94 -225 134 -224
rect 851 -234 891 -233
rect 851 -237 891 -236
rect -148 -283 -147 -243
rect -145 -283 -144 -243
rect -99 -283 -98 -243
rect -96 -283 -95 -243
rect 23 -246 63 -245
rect 23 -249 63 -248
rect 23 -254 63 -253
rect 174 -246 214 -245
rect 851 -242 891 -241
rect 851 -245 891 -244
rect 174 -249 214 -248
rect 23 -257 63 -256
rect -67 -297 -66 -257
rect -64 -297 -63 -257
rect 174 -254 214 -253
rect 396 -253 436 -252
rect 396 -256 436 -255
rect 174 -257 214 -256
rect 396 -261 436 -260
rect 396 -264 436 -263
rect 396 -269 436 -268
rect 780 -266 820 -265
rect 780 -269 820 -268
rect 396 -272 436 -271
rect 94 -278 134 -277
rect 396 -277 436 -276
rect 780 -274 820 -273
rect 931 -266 971 -265
rect 931 -269 971 -268
rect 780 -277 820 -276
rect 396 -280 436 -279
rect 94 -281 134 -280
rect 94 -286 134 -285
rect 931 -274 971 -273
rect 931 -277 971 -276
rect 94 -289 134 -288
rect 851 -298 891 -297
rect 1136 -296 1137 -216
rect 1139 -296 1140 -216
rect 1144 -296 1145 -216
rect 1147 -296 1148 -216
rect 1152 -296 1153 -216
rect 1175 -283 1176 -243
rect 1178 -283 1179 -243
rect 1224 -283 1225 -243
rect 1227 -283 1228 -243
rect 851 -301 891 -300
rect 397 -307 437 -306
rect 851 -306 891 -305
rect 1256 -297 1257 -257
rect 1259 -297 1260 -257
rect 851 -309 891 -308
rect 397 -310 437 -309
rect 94 -316 134 -315
rect 397 -315 437 -314
rect 576 -314 616 -313
rect 576 -317 616 -316
rect 397 -318 437 -317
rect 94 -319 134 -318
rect 94 -324 134 -323
rect 397 -323 437 -322
rect 576 -322 616 -321
rect 576 -325 616 -324
rect 397 -326 437 -325
rect 94 -327 134 -326
rect 576 -330 616 -329
rect 576 -333 616 -332
rect 220 -341 260 -340
rect 576 -338 616 -337
rect 576 -341 616 -340
rect 220 -344 260 -343
rect 851 -345 891 -344
rect 851 -348 891 -347
rect 94 -363 134 -362
rect 396 -356 436 -355
rect 851 -353 891 -352
rect 851 -356 891 -355
rect 396 -359 436 -358
rect 94 -366 134 -365
rect 94 -371 134 -370
rect 396 -364 436 -363
rect 396 -367 436 -366
rect 94 -374 134 -373
rect 780 -377 820 -376
rect 780 -380 820 -379
rect 780 -385 820 -384
rect 931 -377 971 -376
rect 931 -380 971 -379
rect 780 -388 820 -387
rect -387 -486 -386 -406
rect -384 -486 -383 -406
rect -379 -486 -378 -406
rect -376 -486 -375 -406
rect -371 -486 -370 -406
rect 23 -395 63 -394
rect 23 -398 63 -397
rect 23 -403 63 -402
rect 174 -395 214 -394
rect 931 -385 971 -384
rect 931 -388 971 -387
rect 174 -398 214 -397
rect 23 -406 63 -405
rect -348 -473 -347 -433
rect -345 -473 -344 -433
rect -299 -473 -298 -433
rect -296 -473 -295 -433
rect -267 -487 -266 -447
rect -264 -487 -263 -447
rect -186 -487 -185 -407
rect -183 -487 -182 -407
rect -178 -487 -177 -407
rect -175 -487 -174 -407
rect -170 -487 -169 -407
rect 174 -403 214 -402
rect 174 -406 214 -405
rect 851 -409 891 -408
rect 851 -412 891 -411
rect 851 -417 891 -416
rect 851 -420 891 -419
rect 94 -427 134 -426
rect 94 -430 134 -429
rect -147 -474 -146 -434
rect -144 -474 -143 -434
rect -98 -474 -97 -434
rect -95 -474 -94 -434
rect 94 -435 134 -434
rect 396 -427 436 -426
rect 396 -430 436 -429
rect 94 -438 134 -437
rect 396 -435 436 -434
rect 396 -438 436 -437
rect 396 -443 436 -442
rect 396 -446 436 -445
rect -66 -488 -65 -448
rect -63 -488 -62 -448
rect 396 -451 436 -450
rect 396 -454 436 -453
rect 94 -465 134 -464
rect 396 -459 436 -458
rect 396 -462 436 -461
rect 94 -468 134 -467
rect 94 -473 134 -472
rect 94 -476 134 -475
rect 220 -490 260 -489
rect 220 -493 260 -492
rect 396 -490 436 -489
rect 1137 -487 1138 -407
rect 1140 -487 1141 -407
rect 1145 -487 1146 -407
rect 1148 -487 1149 -407
rect 1153 -487 1154 -407
rect 1176 -474 1177 -434
rect 1179 -474 1180 -434
rect 1225 -474 1226 -434
rect 1228 -474 1229 -434
rect 396 -493 436 -492
rect 396 -498 436 -497
rect 396 -501 436 -500
rect 94 -513 134 -512
rect 396 -506 436 -505
rect 1257 -488 1258 -448
rect 1260 -488 1261 -448
rect 396 -509 436 -508
rect 94 -516 134 -515
rect 94 -521 134 -520
rect 396 -514 436 -513
rect 396 -517 436 -516
rect 94 -524 134 -523
rect 23 -545 63 -544
rect 23 -548 63 -547
rect 23 -553 63 -552
rect 174 -545 214 -544
rect 397 -544 437 -543
rect 397 -547 437 -546
rect 174 -548 214 -547
rect 23 -556 63 -555
rect 174 -553 214 -552
rect 397 -552 437 -551
rect 397 -555 437 -554
rect 174 -556 214 -555
rect 397 -560 437 -559
rect 397 -563 437 -562
rect 552 -562 592 -561
rect 552 -565 592 -564
rect 94 -577 134 -576
rect 552 -570 592 -569
rect 552 -573 592 -572
rect 94 -580 134 -579
rect -385 -676 -384 -596
rect -382 -676 -381 -596
rect -377 -676 -376 -596
rect -374 -676 -373 -596
rect -369 -676 -368 -596
rect 94 -585 134 -584
rect 552 -578 592 -577
rect 552 -581 592 -580
rect 94 -588 134 -587
rect 396 -593 436 -592
rect 552 -586 592 -585
rect 552 -589 592 -588
rect 396 -596 436 -595
rect -346 -663 -345 -623
rect -343 -663 -342 -623
rect -297 -663 -296 -623
rect -294 -663 -293 -623
rect -265 -677 -264 -637
rect -262 -677 -261 -637
rect -184 -677 -183 -597
rect -181 -677 -180 -597
rect -176 -677 -175 -597
rect -173 -677 -172 -597
rect -168 -677 -167 -597
rect 396 -601 436 -600
rect 552 -594 592 -593
rect 552 -597 592 -596
rect 396 -604 436 -603
rect 94 -615 134 -614
rect 94 -618 134 -617
rect -145 -664 -144 -624
rect -142 -664 -141 -624
rect -96 -664 -95 -624
rect -93 -664 -92 -624
rect 94 -623 134 -622
rect 94 -626 134 -625
rect -64 -678 -63 -638
rect -61 -678 -60 -638
rect 220 -640 260 -639
rect 220 -643 260 -642
rect 1139 -677 1140 -597
rect 1142 -677 1143 -597
rect 1147 -677 1148 -597
rect 1150 -677 1151 -597
rect 1155 -677 1156 -597
rect 1178 -664 1179 -624
rect 1181 -664 1182 -624
rect 1227 -664 1228 -624
rect 1230 -664 1231 -624
rect 1259 -678 1260 -638
rect 1262 -678 1263 -638
<< ndcontact >>
rect -391 30 -387 50
rect -383 30 -379 50
rect -352 44 -348 84
rect -344 44 -340 84
rect -336 44 -332 84
rect -303 44 -299 84
rect -295 44 -291 84
rect -287 44 -283 84
rect -271 51 -267 71
rect -263 51 -259 71
rect -190 29 -186 49
rect -182 29 -178 49
rect -151 43 -147 83
rect -143 43 -139 83
rect -135 43 -131 83
rect -102 43 -98 83
rect -94 43 -90 83
rect -86 43 -82 83
rect 156 86 196 90
rect 156 78 196 82
rect 156 70 196 74
rect -70 50 -66 70
rect -62 50 -58 70
rect 85 54 125 58
rect 236 54 276 58
rect 85 46 125 50
rect 236 46 276 50
rect 85 38 125 42
rect 236 38 276 42
rect 389 29 393 49
rect 397 29 401 49
rect 428 43 432 83
rect 436 43 440 83
rect 444 43 448 83
rect 477 43 481 83
rect 485 43 489 83
rect 493 43 497 83
rect 509 50 513 70
rect 517 50 521 70
rect 1133 29 1137 49
rect 1141 29 1145 49
rect 1172 43 1176 83
rect 1180 43 1184 83
rect 1188 43 1192 83
rect 1221 43 1225 83
rect 1229 43 1233 83
rect 1237 43 1241 83
rect 1253 50 1257 70
rect 1261 50 1265 70
rect 156 22 196 26
rect 156 14 196 18
rect 156 6 196 10
rect 156 -16 196 -12
rect 913 -14 953 -10
rect 156 -24 196 -20
rect 913 -22 953 -18
rect 156 -32 196 -28
rect 913 -30 953 -26
rect 275 -41 295 -37
rect 458 -40 498 -36
rect 275 -49 295 -45
rect 458 -48 498 -44
rect 625 -48 665 -44
rect 842 -46 882 -42
rect 458 -56 498 -52
rect 156 -63 196 -59
rect 625 -56 665 -52
rect 993 -46 1033 -42
rect 842 -54 882 -50
rect 625 -64 665 -60
rect 993 -54 1033 -50
rect 842 -62 882 -58
rect 993 -62 1033 -58
rect -390 -163 -386 -143
rect -382 -163 -378 -143
rect -351 -149 -347 -109
rect -343 -149 -339 -109
rect -335 -149 -331 -109
rect -302 -149 -298 -109
rect -294 -149 -290 -109
rect -286 -149 -282 -109
rect 156 -71 196 -67
rect 156 -79 196 -75
rect 913 -78 953 -74
rect 913 -86 953 -82
rect 85 -95 125 -91
rect 236 -95 276 -91
rect 913 -94 953 -90
rect 85 -103 125 -99
rect -270 -142 -266 -122
rect -262 -142 -258 -122
rect -189 -164 -185 -144
rect -181 -164 -177 -144
rect -150 -150 -146 -110
rect -142 -150 -138 -110
rect -134 -150 -130 -110
rect -101 -150 -97 -110
rect -93 -150 -89 -110
rect -85 -150 -81 -110
rect 236 -103 276 -99
rect 85 -111 125 -107
rect 236 -111 276 -107
rect -69 -143 -65 -123
rect -61 -143 -57 -123
rect 156 -127 196 -123
rect 913 -123 953 -119
rect 156 -135 196 -131
rect 453 -135 513 -131
rect 913 -131 953 -127
rect 156 -143 196 -139
rect 913 -139 953 -135
rect 453 -143 513 -139
rect 453 -151 513 -147
rect 642 -151 702 -147
rect 453 -159 513 -155
rect 156 -165 196 -161
rect 642 -159 702 -155
rect 842 -155 882 -151
rect 156 -173 196 -169
rect 642 -167 702 -163
rect 993 -155 1033 -151
rect 842 -163 882 -159
rect 993 -163 1033 -159
rect 1134 -164 1138 -144
rect 1142 -164 1146 -144
rect 1173 -150 1177 -110
rect 1181 -150 1185 -110
rect 1189 -150 1193 -110
rect 1222 -150 1226 -110
rect 1230 -150 1234 -110
rect 1238 -150 1242 -110
rect 1254 -143 1258 -123
rect 1262 -143 1266 -123
rect 842 -171 882 -167
rect 993 -171 1033 -167
rect 642 -175 702 -171
rect 156 -181 196 -177
rect 275 -190 295 -186
rect 458 -184 498 -180
rect 275 -198 295 -194
rect 458 -192 498 -188
rect 913 -187 953 -183
rect 458 -200 498 -196
rect 913 -195 953 -191
rect 913 -203 953 -199
rect 156 -213 196 -209
rect 156 -221 196 -217
rect 156 -229 196 -225
rect 913 -233 953 -229
rect 85 -245 125 -241
rect 236 -245 276 -241
rect 913 -241 953 -237
rect 85 -253 125 -249
rect -392 -351 -388 -331
rect -384 -351 -380 -331
rect -353 -337 -349 -297
rect -345 -337 -341 -297
rect -337 -337 -333 -297
rect -304 -337 -300 -297
rect -296 -337 -292 -297
rect -288 -337 -284 -297
rect 236 -253 276 -249
rect 452 -252 532 -248
rect 913 -249 953 -245
rect 85 -261 125 -257
rect 236 -261 276 -257
rect 452 -260 532 -256
rect 452 -268 532 -264
rect 842 -265 882 -261
rect 156 -277 196 -273
rect 452 -276 532 -272
rect 993 -265 1033 -261
rect 842 -273 882 -269
rect 156 -285 196 -281
rect 452 -284 532 -280
rect 993 -273 1033 -269
rect 842 -281 882 -277
rect 993 -281 1033 -277
rect 156 -293 196 -289
rect -272 -330 -268 -310
rect -264 -330 -260 -310
rect -191 -352 -187 -332
rect -183 -352 -179 -332
rect -152 -338 -148 -298
rect -144 -338 -140 -298
rect -136 -338 -132 -298
rect -103 -338 -99 -298
rect -95 -338 -91 -298
rect -87 -338 -83 -298
rect 913 -297 953 -293
rect 453 -306 513 -302
rect 913 -305 953 -301
rect -71 -331 -67 -311
rect -63 -331 -59 -311
rect 156 -315 196 -311
rect 453 -314 513 -310
rect 632 -313 712 -309
rect 913 -313 953 -309
rect 156 -323 196 -319
rect 453 -322 513 -318
rect 632 -321 712 -317
rect 156 -331 196 -327
rect 453 -330 513 -326
rect 632 -329 712 -325
rect 274 -340 294 -336
rect 632 -337 712 -333
rect 274 -348 294 -344
rect 632 -345 712 -341
rect 913 -344 953 -340
rect 156 -362 196 -358
rect 458 -355 498 -351
rect 913 -352 953 -348
rect 1132 -352 1136 -332
rect 1140 -352 1144 -332
rect 1171 -338 1175 -298
rect 1179 -338 1183 -298
rect 1187 -338 1191 -298
rect 1220 -338 1224 -298
rect 1228 -338 1232 -298
rect 1236 -338 1240 -298
rect 1252 -331 1256 -311
rect 1260 -331 1264 -311
rect 156 -370 196 -366
rect 458 -363 498 -359
rect 913 -360 953 -356
rect 458 -371 498 -367
rect 156 -378 196 -374
rect 842 -376 882 -372
rect 993 -376 1033 -372
rect 842 -384 882 -380
rect 85 -394 125 -390
rect 236 -394 276 -390
rect 993 -384 1033 -380
rect 842 -392 882 -388
rect 993 -392 1033 -388
rect 85 -402 125 -398
rect 236 -402 276 -398
rect 85 -410 125 -406
rect 236 -410 276 -406
rect 913 -408 953 -404
rect 913 -416 953 -412
rect 156 -426 196 -422
rect 452 -426 552 -422
rect 913 -424 953 -420
rect 156 -434 196 -430
rect 452 -434 552 -430
rect 156 -442 196 -438
rect 452 -442 552 -438
rect -391 -542 -387 -522
rect -383 -542 -379 -522
rect -352 -528 -348 -488
rect -344 -528 -340 -488
rect -336 -528 -332 -488
rect -303 -528 -299 -488
rect -295 -528 -291 -488
rect -287 -528 -283 -488
rect 452 -450 552 -446
rect 156 -464 196 -460
rect 452 -458 552 -454
rect 452 -466 552 -462
rect 156 -472 196 -468
rect 156 -480 196 -476
rect -271 -521 -267 -501
rect -263 -521 -259 -501
rect -190 -543 -186 -523
rect -182 -543 -178 -523
rect -151 -529 -147 -489
rect -143 -529 -139 -489
rect -135 -529 -131 -489
rect -102 -529 -98 -489
rect -94 -529 -90 -489
rect -86 -529 -82 -489
rect 274 -489 294 -485
rect 452 -489 532 -485
rect 274 -497 294 -493
rect 452 -497 532 -493
rect -70 -522 -66 -502
rect -62 -522 -58 -502
rect 156 -512 196 -508
rect 452 -505 532 -501
rect 156 -520 196 -516
rect 452 -513 532 -509
rect 452 -521 532 -517
rect 156 -528 196 -524
rect 85 -544 125 -540
rect 236 -544 276 -540
rect 453 -543 513 -539
rect 1133 -543 1137 -523
rect 1141 -543 1145 -523
rect 1172 -529 1176 -489
rect 1180 -529 1184 -489
rect 1188 -529 1192 -489
rect 1221 -529 1225 -489
rect 1229 -529 1233 -489
rect 1237 -529 1241 -489
rect 1253 -522 1257 -502
rect 1261 -522 1265 -502
rect 85 -552 125 -548
rect 236 -552 276 -548
rect 453 -551 513 -547
rect 85 -560 125 -556
rect 236 -560 276 -556
rect 453 -559 513 -555
rect 453 -567 513 -563
rect 608 -561 708 -557
rect 156 -576 196 -572
rect 608 -569 708 -565
rect 156 -584 196 -580
rect 608 -577 708 -573
rect 156 -592 196 -588
rect 458 -592 498 -588
rect 608 -585 708 -581
rect 458 -600 498 -596
rect 608 -593 708 -589
rect 608 -601 708 -597
rect 458 -608 498 -604
rect 156 -614 196 -610
rect 156 -622 196 -618
rect 156 -630 196 -626
rect -389 -732 -385 -712
rect -381 -732 -377 -712
rect -350 -718 -346 -678
rect -342 -718 -338 -678
rect -334 -718 -330 -678
rect -301 -718 -297 -678
rect -293 -718 -289 -678
rect -285 -718 -281 -678
rect 274 -639 294 -635
rect 274 -647 294 -643
rect -269 -711 -265 -691
rect -261 -711 -257 -691
rect -188 -733 -184 -713
rect -180 -733 -176 -713
rect -149 -719 -145 -679
rect -141 -719 -137 -679
rect -133 -719 -129 -679
rect -100 -719 -96 -679
rect -92 -719 -88 -679
rect -84 -719 -80 -679
rect -68 -712 -64 -692
rect -60 -712 -56 -692
rect 1135 -733 1139 -713
rect 1143 -733 1147 -713
rect 1174 -719 1178 -679
rect 1182 -719 1186 -679
rect 1190 -719 1194 -679
rect 1223 -719 1227 -679
rect 1231 -719 1235 -679
rect 1239 -719 1243 -679
rect 1255 -712 1259 -692
rect 1263 -712 1267 -692
<< pdcontact >>
rect -391 86 -387 166
rect -383 86 -379 166
rect -375 86 -371 166
rect -352 99 -348 139
rect -344 99 -340 139
rect -303 99 -299 139
rect -295 99 -291 139
rect -271 85 -267 125
rect -263 85 -259 125
rect -190 85 -186 165
rect -182 85 -178 165
rect -174 85 -170 165
rect -151 98 -147 138
rect -143 98 -139 138
rect -102 98 -98 138
rect -94 98 -90 138
rect -70 84 -66 124
rect -62 84 -58 124
rect 94 86 134 90
rect 389 85 393 165
rect 397 85 401 165
rect 405 85 409 165
rect 428 98 432 138
rect 436 98 440 138
rect 477 98 481 138
rect 485 98 489 138
rect 94 78 134 82
rect 94 70 134 74
rect 509 84 513 124
rect 517 84 521 124
rect 1133 85 1137 165
rect 1141 85 1145 165
rect 1149 85 1153 165
rect 1172 98 1176 138
rect 1180 98 1184 138
rect 1221 98 1225 138
rect 1229 98 1233 138
rect 23 54 63 58
rect 174 54 214 58
rect 23 46 63 50
rect 174 46 214 50
rect 23 38 63 42
rect 174 38 214 42
rect 1253 84 1257 124
rect 1261 84 1265 124
rect 94 22 134 26
rect 94 14 134 18
rect 94 6 134 10
rect -390 -107 -386 -27
rect -382 -107 -378 -27
rect -374 -107 -370 -27
rect 94 -16 134 -12
rect 851 -14 891 -10
rect 94 -24 134 -20
rect 851 -22 891 -18
rect -351 -94 -347 -54
rect -343 -94 -339 -54
rect -302 -94 -298 -54
rect -294 -94 -290 -54
rect -270 -108 -266 -68
rect -262 -108 -258 -68
rect -189 -108 -185 -28
rect -181 -108 -177 -28
rect -173 -108 -169 -28
rect 94 -32 134 -28
rect 851 -30 891 -26
rect 221 -41 261 -37
rect 396 -40 436 -36
rect 221 -49 261 -45
rect 396 -48 436 -44
rect 563 -48 603 -44
rect -150 -95 -146 -55
rect -142 -95 -138 -55
rect -101 -95 -97 -55
rect -93 -95 -89 -55
rect 396 -56 436 -52
rect 780 -46 820 -42
rect 931 -46 971 -42
rect 563 -56 603 -52
rect 94 -63 134 -59
rect 780 -54 820 -50
rect 931 -54 971 -50
rect 563 -64 603 -60
rect 780 -62 820 -58
rect 931 -62 971 -58
rect -69 -109 -65 -69
rect -61 -109 -57 -69
rect 94 -71 134 -67
rect 94 -79 134 -75
rect 851 -78 891 -74
rect 851 -86 891 -82
rect 23 -95 63 -91
rect 174 -95 214 -91
rect 23 -103 63 -99
rect 851 -94 891 -90
rect 174 -103 214 -99
rect 23 -111 63 -107
rect 174 -111 214 -107
rect 1134 -108 1138 -28
rect 1142 -108 1146 -28
rect 1150 -108 1154 -28
rect 1173 -95 1177 -55
rect 1181 -95 1185 -55
rect 1222 -95 1226 -55
rect 1230 -95 1234 -55
rect 1254 -109 1258 -69
rect 1262 -109 1266 -69
rect 851 -123 891 -119
rect 94 -127 134 -123
rect 94 -135 134 -131
rect 851 -131 891 -127
rect 397 -135 437 -131
rect 94 -143 134 -139
rect 397 -143 437 -139
rect 851 -139 891 -135
rect 397 -151 437 -147
rect 586 -151 626 -147
rect 397 -159 437 -155
rect 586 -159 626 -155
rect 94 -165 134 -161
rect 780 -155 820 -151
rect 931 -155 971 -151
rect 586 -167 626 -163
rect 94 -173 134 -169
rect 780 -163 820 -159
rect 931 -163 971 -159
rect 586 -175 626 -171
rect 780 -171 820 -167
rect 931 -171 971 -167
rect 94 -181 134 -177
rect 396 -184 436 -180
rect 221 -190 261 -186
rect 851 -187 891 -183
rect 396 -192 436 -188
rect 221 -198 261 -194
rect 851 -195 891 -191
rect 396 -200 436 -196
rect 851 -203 891 -199
rect -392 -295 -388 -215
rect -384 -295 -380 -215
rect -376 -295 -372 -215
rect 94 -213 134 -209
rect -353 -282 -349 -242
rect -345 -282 -341 -242
rect -304 -282 -300 -242
rect -296 -282 -292 -242
rect -272 -296 -268 -256
rect -264 -296 -260 -256
rect -191 -296 -187 -216
rect -183 -296 -179 -216
rect -175 -296 -171 -216
rect 94 -221 134 -217
rect 94 -229 134 -225
rect 851 -233 891 -229
rect 851 -241 891 -237
rect -152 -283 -148 -243
rect -144 -283 -140 -243
rect -103 -283 -99 -243
rect -95 -283 -91 -243
rect 23 -245 63 -241
rect 174 -245 214 -241
rect 23 -253 63 -249
rect 174 -253 214 -249
rect -71 -297 -67 -257
rect -63 -297 -59 -257
rect 23 -261 63 -257
rect 396 -252 436 -248
rect 851 -249 891 -245
rect 174 -261 214 -257
rect 396 -260 436 -256
rect 396 -268 436 -264
rect 780 -265 820 -261
rect 931 -265 971 -261
rect 94 -277 134 -273
rect 396 -276 436 -272
rect 780 -273 820 -269
rect 931 -273 971 -269
rect 94 -285 134 -281
rect 396 -284 436 -280
rect 780 -281 820 -277
rect 931 -281 971 -277
rect 94 -293 134 -289
rect 851 -297 891 -293
rect 1132 -296 1136 -216
rect 1140 -296 1144 -216
rect 1148 -296 1152 -216
rect 1171 -283 1175 -243
rect 1179 -283 1183 -243
rect 1220 -283 1224 -243
rect 1228 -283 1232 -243
rect 397 -306 437 -302
rect 851 -305 891 -301
rect 1252 -297 1256 -257
rect 1260 -297 1264 -257
rect 94 -315 134 -311
rect 397 -314 437 -310
rect 576 -313 616 -309
rect 851 -313 891 -309
rect 94 -323 134 -319
rect 397 -322 437 -318
rect 576 -321 616 -317
rect 94 -331 134 -327
rect 397 -330 437 -326
rect 576 -329 616 -325
rect 220 -340 260 -336
rect 576 -337 616 -333
rect 220 -348 260 -344
rect 576 -345 616 -341
rect 851 -344 891 -340
rect 396 -355 436 -351
rect 94 -362 134 -358
rect 851 -352 891 -348
rect 396 -363 436 -359
rect 94 -370 134 -366
rect 851 -360 891 -356
rect 396 -371 436 -367
rect 94 -378 134 -374
rect 780 -376 820 -372
rect 931 -376 971 -372
rect 780 -384 820 -380
rect 931 -384 971 -380
rect 23 -394 63 -390
rect -391 -486 -387 -406
rect -383 -486 -379 -406
rect -375 -486 -371 -406
rect 174 -394 214 -390
rect 23 -402 63 -398
rect 780 -392 820 -388
rect 931 -392 971 -388
rect 174 -402 214 -398
rect -352 -473 -348 -433
rect -344 -473 -340 -433
rect -303 -473 -299 -433
rect -295 -473 -291 -433
rect -271 -487 -267 -447
rect -263 -487 -259 -447
rect -190 -487 -186 -407
rect -182 -487 -178 -407
rect -174 -487 -170 -407
rect 23 -410 63 -406
rect 174 -410 214 -406
rect 851 -408 891 -404
rect 851 -416 891 -412
rect 94 -426 134 -422
rect 396 -426 436 -422
rect 94 -434 134 -430
rect -151 -474 -147 -434
rect -143 -474 -139 -434
rect -102 -474 -98 -434
rect -94 -474 -90 -434
rect 851 -424 891 -420
rect 396 -434 436 -430
rect 94 -442 134 -438
rect 396 -442 436 -438
rect -70 -488 -66 -448
rect -62 -488 -58 -448
rect 396 -450 436 -446
rect 396 -458 436 -454
rect 94 -464 134 -460
rect 396 -466 436 -462
rect 94 -472 134 -468
rect 94 -480 134 -476
rect 220 -489 260 -485
rect 396 -489 436 -485
rect 220 -497 260 -493
rect 1133 -487 1137 -407
rect 1141 -487 1145 -407
rect 1149 -487 1153 -407
rect 1172 -474 1176 -434
rect 1180 -474 1184 -434
rect 1221 -474 1225 -434
rect 1229 -474 1233 -434
rect 396 -497 436 -493
rect 396 -505 436 -501
rect 94 -512 134 -508
rect 1253 -488 1257 -448
rect 1261 -488 1265 -448
rect 396 -513 436 -509
rect 94 -520 134 -516
rect 396 -521 436 -517
rect 94 -528 134 -524
rect 23 -544 63 -540
rect 174 -544 214 -540
rect 23 -552 63 -548
rect 397 -543 437 -539
rect 174 -552 214 -548
rect 23 -560 63 -556
rect 397 -551 437 -547
rect 174 -560 214 -556
rect 397 -559 437 -555
rect 552 -561 592 -557
rect 397 -567 437 -563
rect 552 -569 592 -565
rect 94 -576 134 -572
rect 552 -577 592 -573
rect 94 -584 134 -580
rect -389 -676 -385 -596
rect -381 -676 -377 -596
rect -373 -676 -369 -596
rect 552 -585 592 -581
rect 94 -592 134 -588
rect 396 -592 436 -588
rect 552 -593 592 -589
rect -350 -663 -346 -623
rect -342 -663 -338 -623
rect -301 -663 -297 -623
rect -293 -663 -289 -623
rect -269 -677 -265 -637
rect -261 -677 -257 -637
rect -188 -677 -184 -597
rect -180 -677 -176 -597
rect -172 -677 -168 -597
rect 396 -600 436 -596
rect 552 -601 592 -597
rect 396 -608 436 -604
rect 94 -614 134 -610
rect 94 -622 134 -618
rect -149 -664 -145 -624
rect -141 -664 -137 -624
rect -100 -664 -96 -624
rect -92 -664 -88 -624
rect 94 -630 134 -626
rect -68 -678 -64 -638
rect -60 -678 -56 -638
rect 220 -639 260 -635
rect 220 -647 260 -643
rect 1135 -677 1139 -597
rect 1143 -677 1147 -597
rect 1151 -677 1155 -597
rect 1174 -664 1178 -624
rect 1182 -664 1186 -624
rect 1223 -664 1227 -624
rect 1231 -664 1235 -624
rect 1255 -678 1259 -638
rect 1263 -678 1267 -638
<< polysilicon >>
rect -386 166 -384 172
rect -378 166 -376 179
rect -185 165 -183 171
rect -177 165 -175 178
rect 394 165 396 171
rect 402 165 404 178
rect 1138 165 1140 171
rect 1146 165 1148 178
rect -347 139 -345 150
rect -298 139 -296 150
rect -266 125 -264 128
rect -386 79 -384 86
rect -385 75 -384 79
rect -378 75 -376 86
rect -347 84 -345 99
rect -339 84 -337 87
rect -298 84 -296 99
rect -290 84 -288 87
rect -146 138 -144 149
rect -97 138 -95 149
rect -65 124 -63 127
rect -386 50 -384 75
rect -266 71 -264 85
rect -185 78 -183 85
rect -184 74 -183 78
rect -177 74 -175 85
rect -146 83 -144 98
rect -138 83 -136 86
rect -97 83 -95 98
rect -89 83 -87 86
rect -266 48 -264 51
rect -185 49 -183 74
rect -347 40 -345 44
rect -339 40 -337 44
rect -298 40 -296 44
rect -290 40 -288 44
rect -386 26 -384 30
rect -65 70 -63 84
rect 433 138 435 149
rect 482 138 484 149
rect 514 124 516 127
rect 81 83 94 85
rect 134 83 156 85
rect 196 83 199 85
rect 394 78 396 85
rect 81 75 94 77
rect 134 75 156 77
rect 196 75 199 77
rect 395 74 396 78
rect 402 74 404 85
rect 433 83 435 98
rect 441 83 443 86
rect 482 83 484 98
rect 490 83 492 86
rect 1177 138 1179 149
rect 1226 138 1228 149
rect 1258 124 1260 127
rect 10 51 23 53
rect 63 51 85 53
rect 125 51 128 53
rect -65 47 -63 50
rect -146 39 -144 43
rect -138 39 -136 43
rect -97 39 -95 43
rect -89 39 -87 43
rect 161 51 174 53
rect 214 51 236 53
rect 276 51 279 53
rect 10 43 23 45
rect 63 43 85 45
rect 125 43 128 45
rect 394 49 396 74
rect 161 43 174 45
rect 214 43 236 45
rect 276 43 279 45
rect 514 70 516 84
rect 1138 78 1140 85
rect 1139 74 1140 78
rect 1146 74 1148 85
rect 1177 83 1179 98
rect 1185 83 1187 86
rect 1226 83 1228 98
rect 1234 83 1236 86
rect 514 47 516 50
rect 1138 49 1140 74
rect 433 39 435 43
rect 441 39 443 43
rect 482 39 484 43
rect 490 39 492 43
rect 1258 70 1260 84
rect 1258 47 1260 50
rect 1177 39 1179 43
rect 1185 39 1187 43
rect 1226 39 1228 43
rect 1234 39 1236 43
rect -185 25 -183 29
rect 394 25 396 29
rect 1138 25 1140 29
rect 81 19 94 21
rect 134 19 156 21
rect 196 19 199 21
rect 81 11 94 13
rect 134 11 156 13
rect 196 11 199 13
rect -385 -27 -383 -21
rect -377 -27 -375 -14
rect -184 -28 -182 -22
rect -176 -28 -174 -15
rect 81 -19 94 -17
rect 134 -19 156 -17
rect 196 -19 199 -17
rect 838 -17 851 -15
rect 891 -17 913 -15
rect 953 -17 956 -15
rect 81 -27 94 -25
rect 134 -27 156 -25
rect 196 -27 199 -25
rect 838 -25 851 -23
rect 891 -25 913 -23
rect 953 -25 956 -23
rect -346 -54 -344 -43
rect -297 -54 -295 -43
rect -265 -68 -263 -65
rect -385 -114 -383 -107
rect -384 -118 -383 -114
rect -377 -118 -375 -107
rect -346 -109 -344 -94
rect -338 -109 -336 -106
rect -297 -109 -295 -94
rect -289 -109 -287 -106
rect 1139 -28 1141 -22
rect 1147 -28 1149 -15
rect 201 -44 221 -42
rect 261 -44 275 -42
rect 295 -44 298 -42
rect 383 -43 396 -41
rect 436 -43 458 -41
rect 498 -43 501 -41
rect -145 -55 -143 -44
rect -96 -55 -94 -44
rect 383 -51 396 -49
rect 436 -51 458 -49
rect 498 -51 501 -49
rect 550 -51 563 -49
rect 603 -51 625 -49
rect 665 -51 668 -49
rect 767 -49 780 -47
rect 820 -49 842 -47
rect 882 -49 885 -47
rect -64 -69 -62 -66
rect 550 -59 563 -57
rect 603 -59 625 -57
rect 665 -59 668 -57
rect 918 -49 931 -47
rect 971 -49 993 -47
rect 1033 -49 1036 -47
rect 767 -57 780 -55
rect 820 -57 842 -55
rect 882 -57 885 -55
rect 918 -57 931 -55
rect 971 -57 993 -55
rect 1033 -57 1036 -55
rect 81 -66 94 -64
rect 134 -66 156 -64
rect 196 -66 199 -64
rect -385 -143 -383 -118
rect -265 -122 -263 -108
rect -184 -115 -182 -108
rect -183 -119 -182 -115
rect -176 -119 -174 -108
rect -145 -110 -143 -95
rect -137 -110 -135 -107
rect -96 -110 -94 -95
rect -88 -110 -86 -107
rect 81 -74 94 -72
rect 134 -74 156 -72
rect 196 -74 199 -72
rect 838 -81 851 -79
rect 891 -81 913 -79
rect 953 -81 956 -79
rect 838 -89 851 -87
rect 891 -89 913 -87
rect 953 -89 956 -87
rect 10 -98 23 -96
rect 63 -98 85 -96
rect 125 -98 128 -96
rect 161 -98 174 -96
rect 214 -98 236 -96
rect 276 -98 279 -96
rect 10 -106 23 -104
rect 63 -106 85 -104
rect 125 -106 128 -104
rect -265 -145 -263 -142
rect -184 -144 -182 -119
rect -346 -153 -344 -149
rect -338 -153 -336 -149
rect -297 -153 -295 -149
rect -289 -153 -287 -149
rect -385 -167 -383 -163
rect -64 -123 -62 -109
rect 161 -106 174 -104
rect 214 -106 236 -104
rect 276 -106 279 -104
rect 1178 -55 1180 -44
rect 1227 -55 1229 -44
rect 1259 -69 1261 -66
rect 1139 -115 1141 -108
rect 1140 -119 1141 -115
rect 1147 -119 1149 -108
rect 1178 -110 1180 -95
rect 1186 -110 1188 -107
rect 1227 -110 1229 -95
rect 1235 -110 1237 -107
rect 838 -126 851 -124
rect 891 -126 913 -124
rect 953 -126 956 -124
rect 81 -130 94 -128
rect 134 -130 156 -128
rect 196 -130 199 -128
rect 81 -138 94 -136
rect 134 -138 156 -136
rect 196 -138 199 -136
rect 838 -134 851 -132
rect 891 -134 913 -132
rect 953 -134 956 -132
rect 383 -138 397 -136
rect 437 -138 453 -136
rect 513 -138 516 -136
rect -64 -146 -62 -143
rect 1139 -144 1141 -119
rect 383 -146 397 -144
rect 437 -146 453 -144
rect 513 -146 516 -144
rect -145 -154 -143 -150
rect -137 -154 -135 -150
rect -96 -154 -94 -150
rect -88 -154 -86 -150
rect 383 -154 397 -152
rect 437 -154 453 -152
rect 513 -154 516 -152
rect 572 -154 586 -152
rect 626 -154 642 -152
rect 702 -154 705 -152
rect -184 -168 -182 -164
rect 767 -158 780 -156
rect 820 -158 842 -156
rect 882 -158 885 -156
rect 572 -162 586 -160
rect 626 -162 642 -160
rect 702 -162 705 -160
rect 81 -168 94 -166
rect 134 -168 156 -166
rect 196 -168 199 -166
rect 918 -158 931 -156
rect 971 -158 993 -156
rect 1033 -158 1036 -156
rect 767 -166 780 -164
rect 820 -166 842 -164
rect 882 -166 885 -164
rect 572 -170 586 -168
rect 626 -170 642 -168
rect 702 -170 705 -168
rect 81 -176 94 -174
rect 134 -176 156 -174
rect 196 -176 199 -174
rect 1259 -123 1261 -109
rect 1259 -146 1261 -143
rect 1178 -154 1180 -150
rect 1186 -154 1188 -150
rect 1227 -154 1229 -150
rect 1235 -154 1237 -150
rect 918 -166 931 -164
rect 971 -166 993 -164
rect 1033 -166 1036 -164
rect 1139 -168 1141 -164
rect 383 -187 396 -185
rect 436 -187 458 -185
rect 498 -187 501 -185
rect 201 -193 221 -191
rect 261 -193 275 -191
rect 295 -193 298 -191
rect 838 -190 851 -188
rect 891 -190 913 -188
rect 953 -190 956 -188
rect 383 -195 396 -193
rect 436 -195 458 -193
rect 498 -195 501 -193
rect -387 -215 -385 -209
rect -379 -215 -377 -202
rect 838 -198 851 -196
rect 891 -198 913 -196
rect 953 -198 956 -196
rect -186 -216 -184 -210
rect -178 -216 -176 -203
rect -348 -242 -346 -231
rect -299 -242 -297 -231
rect -267 -256 -265 -253
rect -387 -302 -385 -295
rect -386 -306 -385 -302
rect -379 -306 -377 -295
rect -348 -297 -346 -282
rect -340 -297 -338 -294
rect -299 -297 -297 -282
rect -291 -297 -289 -294
rect 81 -216 94 -214
rect 134 -216 156 -214
rect 196 -216 199 -214
rect 1137 -216 1139 -210
rect 1145 -216 1147 -203
rect 81 -224 94 -222
rect 134 -224 156 -222
rect 196 -224 199 -222
rect -147 -243 -145 -232
rect -98 -243 -96 -232
rect 838 -236 851 -234
rect 891 -236 913 -234
rect 953 -236 956 -234
rect 10 -248 23 -246
rect 63 -248 85 -246
rect 125 -248 128 -246
rect -66 -257 -64 -254
rect 838 -244 851 -242
rect 891 -244 913 -242
rect 953 -244 956 -242
rect 161 -248 174 -246
rect 214 -248 236 -246
rect 276 -248 279 -246
rect 10 -256 23 -254
rect 63 -256 85 -254
rect 125 -256 128 -254
rect -387 -331 -385 -306
rect -267 -310 -265 -296
rect -186 -303 -184 -296
rect -185 -307 -184 -303
rect -178 -307 -176 -296
rect -147 -298 -145 -283
rect -139 -298 -137 -295
rect -98 -298 -96 -283
rect -90 -298 -88 -295
rect 161 -256 174 -254
rect 214 -256 236 -254
rect 276 -256 279 -254
rect 383 -255 396 -253
rect 436 -255 452 -253
rect 532 -255 535 -253
rect 383 -263 396 -261
rect 436 -263 452 -261
rect 532 -263 535 -261
rect 767 -268 780 -266
rect 820 -268 842 -266
rect 882 -268 885 -266
rect 383 -271 396 -269
rect 436 -271 452 -269
rect 532 -271 535 -269
rect 81 -280 94 -278
rect 134 -280 156 -278
rect 196 -280 199 -278
rect 918 -268 931 -266
rect 971 -268 993 -266
rect 1033 -268 1036 -266
rect 767 -276 780 -274
rect 820 -276 842 -274
rect 882 -276 885 -274
rect 383 -279 396 -277
rect 436 -279 452 -277
rect 532 -279 535 -277
rect 918 -276 931 -274
rect 971 -276 993 -274
rect 1033 -276 1036 -274
rect 81 -288 94 -286
rect 134 -288 156 -286
rect 196 -288 199 -286
rect -267 -333 -265 -330
rect -186 -332 -184 -307
rect -348 -341 -346 -337
rect -340 -341 -338 -337
rect -299 -341 -297 -337
rect -291 -341 -289 -337
rect -387 -355 -385 -351
rect -66 -311 -64 -297
rect 1176 -243 1178 -232
rect 1225 -243 1227 -232
rect 1257 -257 1259 -254
rect 838 -300 851 -298
rect 891 -300 913 -298
rect 953 -300 956 -298
rect 383 -309 397 -307
rect 437 -309 453 -307
rect 513 -309 516 -307
rect 1137 -303 1139 -296
rect 838 -308 851 -306
rect 891 -308 913 -306
rect 953 -308 956 -306
rect 1138 -307 1139 -303
rect 1145 -307 1147 -296
rect 1176 -298 1178 -283
rect 1184 -298 1186 -295
rect 1225 -298 1227 -283
rect 1233 -298 1235 -295
rect 81 -318 94 -316
rect 134 -318 156 -316
rect 196 -318 199 -316
rect 383 -317 397 -315
rect 437 -317 453 -315
rect 513 -317 516 -315
rect 563 -316 576 -314
rect 616 -316 632 -314
rect 712 -316 715 -314
rect 81 -326 94 -324
rect 134 -326 156 -324
rect 196 -326 199 -324
rect 383 -325 397 -323
rect 437 -325 453 -323
rect 513 -325 516 -323
rect 563 -324 576 -322
rect 616 -324 632 -322
rect 712 -324 715 -322
rect -66 -334 -64 -331
rect 563 -332 576 -330
rect 616 -332 632 -330
rect 712 -332 715 -330
rect 1137 -332 1139 -307
rect -147 -342 -145 -338
rect -139 -342 -137 -338
rect -98 -342 -96 -338
rect -90 -342 -88 -338
rect 563 -340 576 -338
rect 616 -340 632 -338
rect 712 -340 715 -338
rect 200 -343 220 -341
rect 260 -343 274 -341
rect 294 -343 297 -341
rect 838 -347 851 -345
rect 891 -347 913 -345
rect 953 -347 956 -345
rect -186 -356 -184 -352
rect 1257 -311 1259 -297
rect 1257 -334 1259 -331
rect 1176 -342 1178 -338
rect 1184 -342 1186 -338
rect 1225 -342 1227 -338
rect 1233 -342 1235 -338
rect 838 -355 851 -353
rect 891 -355 913 -353
rect 953 -355 956 -353
rect 383 -358 396 -356
rect 436 -358 458 -356
rect 498 -358 501 -356
rect 81 -365 94 -363
rect 134 -365 156 -363
rect 196 -365 199 -363
rect 1137 -356 1139 -352
rect 383 -366 396 -364
rect 436 -366 458 -364
rect 498 -366 501 -364
rect 81 -373 94 -371
rect 134 -373 156 -371
rect 196 -373 199 -371
rect 767 -379 780 -377
rect 820 -379 842 -377
rect 882 -379 885 -377
rect 918 -379 931 -377
rect 971 -379 993 -377
rect 1033 -379 1036 -377
rect 767 -387 780 -385
rect 820 -387 842 -385
rect 882 -387 885 -385
rect -386 -406 -384 -400
rect -378 -406 -376 -393
rect -185 -407 -183 -401
rect -177 -407 -175 -394
rect 10 -397 23 -395
rect 63 -397 85 -395
rect 125 -397 128 -395
rect 918 -387 931 -385
rect 971 -387 993 -385
rect 1033 -387 1036 -385
rect 161 -397 174 -395
rect 214 -397 236 -395
rect 276 -397 279 -395
rect 10 -405 23 -403
rect 63 -405 85 -403
rect 125 -405 128 -403
rect -347 -433 -345 -422
rect -298 -433 -296 -422
rect -266 -447 -264 -444
rect -386 -493 -384 -486
rect -385 -497 -384 -493
rect -378 -497 -376 -486
rect -347 -488 -345 -473
rect -339 -488 -337 -485
rect -298 -488 -296 -473
rect -290 -488 -288 -485
rect 161 -405 174 -403
rect 214 -405 236 -403
rect 276 -405 279 -403
rect 1138 -407 1140 -401
rect 1146 -407 1148 -394
rect 838 -411 851 -409
rect 891 -411 913 -409
rect 953 -411 956 -409
rect 838 -419 851 -417
rect 891 -419 913 -417
rect 953 -419 956 -417
rect -146 -434 -144 -423
rect -97 -434 -95 -423
rect 81 -429 94 -427
rect 134 -429 156 -427
rect 196 -429 199 -427
rect 383 -429 396 -427
rect 436 -429 452 -427
rect 552 -429 555 -427
rect 81 -437 94 -435
rect 134 -437 156 -435
rect 196 -437 199 -435
rect 383 -437 396 -435
rect 436 -437 452 -435
rect 552 -437 555 -435
rect -65 -448 -63 -445
rect 383 -445 396 -443
rect 436 -445 452 -443
rect 552 -445 555 -443
rect -386 -522 -384 -497
rect -266 -501 -264 -487
rect -185 -494 -183 -487
rect -184 -498 -183 -494
rect -177 -498 -175 -487
rect -146 -489 -144 -474
rect -138 -489 -136 -486
rect -97 -489 -95 -474
rect -89 -489 -87 -486
rect 383 -453 396 -451
rect 436 -453 452 -451
rect 552 -453 555 -451
rect 383 -461 396 -459
rect 436 -461 452 -459
rect 552 -461 555 -459
rect 81 -467 94 -465
rect 134 -467 156 -465
rect 196 -467 199 -465
rect 81 -475 94 -473
rect 134 -475 156 -473
rect 196 -475 199 -473
rect -266 -524 -264 -521
rect -185 -523 -183 -498
rect -347 -532 -345 -528
rect -339 -532 -337 -528
rect -298 -532 -296 -528
rect -290 -532 -288 -528
rect -386 -546 -384 -542
rect -65 -502 -63 -488
rect 200 -492 220 -490
rect 260 -492 274 -490
rect 294 -492 297 -490
rect 1177 -434 1179 -423
rect 1226 -434 1228 -423
rect 1258 -448 1260 -445
rect 383 -492 396 -490
rect 436 -492 452 -490
rect 532 -492 535 -490
rect 1138 -494 1140 -487
rect 383 -500 396 -498
rect 436 -500 452 -498
rect 532 -500 535 -498
rect 1139 -498 1140 -494
rect 1146 -498 1148 -487
rect 1177 -489 1179 -474
rect 1185 -489 1187 -486
rect 1226 -489 1228 -474
rect 1234 -489 1236 -486
rect 383 -508 396 -506
rect 436 -508 452 -506
rect 532 -508 535 -506
rect 81 -515 94 -513
rect 134 -515 156 -513
rect 196 -515 199 -513
rect -65 -525 -63 -522
rect 383 -516 396 -514
rect 436 -516 452 -514
rect 532 -516 535 -514
rect 81 -523 94 -521
rect 134 -523 156 -521
rect 196 -523 199 -521
rect 1138 -523 1140 -498
rect -146 -533 -144 -529
rect -138 -533 -136 -529
rect -97 -533 -95 -529
rect -89 -533 -87 -529
rect -185 -547 -183 -543
rect 10 -547 23 -545
rect 63 -547 85 -545
rect 125 -547 128 -545
rect 161 -547 174 -545
rect 214 -547 236 -545
rect 276 -547 279 -545
rect 1258 -502 1260 -488
rect 1258 -525 1260 -522
rect 1177 -533 1179 -529
rect 1185 -533 1187 -529
rect 1226 -533 1228 -529
rect 1234 -533 1236 -529
rect 383 -546 397 -544
rect 437 -546 453 -544
rect 513 -546 516 -544
rect 10 -555 23 -553
rect 63 -555 85 -553
rect 125 -555 128 -553
rect 161 -555 174 -553
rect 214 -555 236 -553
rect 276 -555 279 -553
rect 1138 -547 1140 -543
rect 383 -554 397 -552
rect 437 -554 453 -552
rect 513 -554 516 -552
rect 383 -562 397 -560
rect 437 -562 453 -560
rect 513 -562 516 -560
rect 539 -564 552 -562
rect 592 -564 608 -562
rect 708 -564 711 -562
rect 539 -572 552 -570
rect 592 -572 608 -570
rect 708 -572 711 -570
rect 81 -579 94 -577
rect 134 -579 156 -577
rect 196 -579 199 -577
rect -384 -596 -382 -590
rect -376 -596 -374 -583
rect -183 -597 -181 -591
rect -175 -597 -173 -584
rect 539 -580 552 -578
rect 592 -580 608 -578
rect 708 -580 711 -578
rect 81 -587 94 -585
rect 134 -587 156 -585
rect 196 -587 199 -585
rect 539 -588 552 -586
rect 592 -588 608 -586
rect 708 -588 711 -586
rect 383 -595 396 -593
rect 436 -595 458 -593
rect 498 -595 501 -593
rect -345 -623 -343 -612
rect -296 -623 -294 -612
rect -264 -637 -262 -634
rect -384 -683 -382 -676
rect -383 -687 -382 -683
rect -376 -687 -374 -676
rect -345 -678 -343 -663
rect -337 -678 -335 -675
rect -296 -678 -294 -663
rect -288 -678 -286 -675
rect 539 -596 552 -594
rect 592 -596 608 -594
rect 708 -596 711 -594
rect 1140 -597 1142 -591
rect 1148 -597 1150 -584
rect 383 -603 396 -601
rect 436 -603 458 -601
rect 498 -603 501 -601
rect -144 -624 -142 -613
rect -95 -624 -93 -613
rect 81 -617 94 -615
rect 134 -617 156 -615
rect 196 -617 199 -615
rect 81 -625 94 -623
rect 134 -625 156 -623
rect 196 -625 199 -623
rect -63 -638 -61 -635
rect -384 -712 -382 -687
rect -264 -691 -262 -677
rect -183 -684 -181 -677
rect -182 -688 -181 -684
rect -175 -688 -173 -677
rect -144 -679 -142 -664
rect -136 -679 -134 -676
rect -95 -679 -93 -664
rect -87 -679 -85 -676
rect 200 -642 220 -640
rect 260 -642 274 -640
rect 294 -642 297 -640
rect 1179 -624 1181 -613
rect 1228 -624 1230 -613
rect 1260 -638 1262 -635
rect -264 -714 -262 -711
rect -183 -713 -181 -688
rect -345 -722 -343 -718
rect -337 -722 -335 -718
rect -296 -722 -294 -718
rect -288 -722 -286 -718
rect -384 -736 -382 -732
rect -63 -692 -61 -678
rect 1140 -684 1142 -677
rect 1141 -688 1142 -684
rect 1148 -688 1150 -677
rect 1179 -679 1181 -664
rect 1187 -679 1189 -676
rect 1228 -679 1230 -664
rect 1236 -679 1238 -676
rect -63 -715 -61 -712
rect 1140 -713 1142 -688
rect -144 -723 -142 -719
rect -136 -723 -134 -719
rect -95 -723 -93 -719
rect -87 -723 -85 -719
rect 1260 -692 1262 -678
rect 1260 -715 1262 -712
rect 1179 -723 1181 -719
rect 1187 -723 1189 -719
rect 1228 -723 1230 -719
rect 1236 -723 1238 -719
rect -183 -737 -181 -733
rect 1140 -737 1142 -733
<< polycontact >>
rect -379 179 -375 183
rect -178 178 -174 182
rect 401 178 405 182
rect 1145 178 1149 182
rect -348 150 -344 154
rect -299 150 -295 154
rect -389 75 -385 79
rect -340 87 -336 91
rect -291 87 -287 91
rect -147 149 -143 153
rect -98 149 -94 153
rect -270 74 -266 78
rect -188 74 -184 78
rect -139 86 -135 90
rect -90 86 -86 90
rect -69 73 -65 77
rect 77 82 81 86
rect 432 149 436 153
rect 481 149 485 153
rect 77 74 81 78
rect 391 74 395 78
rect 440 86 444 90
rect 489 86 493 90
rect 1176 149 1180 153
rect 1225 149 1229 153
rect 6 50 10 54
rect 6 42 10 46
rect 157 50 161 54
rect 157 42 161 46
rect 510 73 514 77
rect 1135 74 1139 78
rect 1184 86 1188 90
rect 1233 86 1237 90
rect 1254 73 1258 77
rect 77 18 81 22
rect 77 10 81 14
rect -378 -14 -374 -10
rect -177 -15 -173 -11
rect 77 -20 81 -16
rect 834 -18 838 -14
rect 1146 -15 1150 -11
rect 77 -28 81 -24
rect 834 -26 838 -22
rect -347 -43 -343 -39
rect -298 -43 -294 -39
rect -388 -118 -384 -114
rect -339 -106 -335 -102
rect -290 -106 -286 -102
rect -146 -44 -142 -40
rect -97 -44 -93 -40
rect 201 -42 205 -38
rect 379 -44 383 -40
rect 379 -52 383 -48
rect 546 -52 550 -48
rect 763 -50 767 -46
rect 77 -67 81 -63
rect 546 -60 550 -56
rect 763 -58 767 -54
rect 914 -50 918 -46
rect 914 -58 918 -54
rect -269 -119 -265 -115
rect -187 -119 -183 -115
rect -138 -107 -134 -103
rect -89 -107 -85 -103
rect 77 -75 81 -71
rect 834 -82 838 -78
rect 834 -90 838 -86
rect 6 -99 10 -95
rect 6 -107 10 -103
rect 157 -99 161 -95
rect -68 -120 -64 -116
rect 157 -107 161 -103
rect 1177 -44 1181 -40
rect 1226 -44 1230 -40
rect 1136 -119 1140 -115
rect 1185 -107 1189 -103
rect 1234 -107 1238 -103
rect 77 -131 81 -127
rect 834 -127 838 -123
rect 77 -139 81 -135
rect 379 -139 383 -135
rect 834 -135 838 -131
rect 379 -147 383 -143
rect 379 -155 383 -151
rect 568 -155 572 -151
rect 77 -169 81 -165
rect 568 -163 572 -159
rect 763 -159 767 -155
rect 77 -177 81 -173
rect 568 -171 572 -167
rect 763 -167 767 -163
rect 914 -159 918 -155
rect 914 -167 918 -163
rect 1255 -120 1259 -116
rect 201 -191 205 -187
rect 379 -188 383 -184
rect 379 -196 383 -192
rect 834 -191 838 -187
rect -380 -202 -376 -198
rect -179 -203 -175 -199
rect 834 -199 838 -195
rect 1144 -203 1148 -199
rect -349 -231 -345 -227
rect -300 -231 -296 -227
rect -390 -306 -386 -302
rect -341 -294 -337 -290
rect -292 -294 -288 -290
rect 77 -217 81 -213
rect 77 -225 81 -221
rect -148 -232 -144 -228
rect -99 -232 -95 -228
rect 834 -237 838 -233
rect 6 -249 10 -245
rect 6 -257 10 -253
rect 157 -249 161 -245
rect 834 -245 838 -241
rect -271 -307 -267 -303
rect -189 -307 -185 -303
rect -140 -295 -136 -291
rect -91 -295 -87 -291
rect 157 -257 161 -253
rect 379 -256 383 -252
rect 379 -264 383 -260
rect 379 -272 383 -268
rect 763 -269 767 -265
rect 77 -281 81 -277
rect 379 -280 383 -276
rect 763 -277 767 -273
rect 914 -269 918 -265
rect 77 -289 81 -285
rect 914 -277 918 -273
rect -70 -308 -66 -304
rect 834 -301 838 -297
rect 1175 -232 1179 -228
rect 1224 -232 1228 -228
rect 379 -310 383 -306
rect 834 -309 838 -305
rect 1134 -307 1138 -303
rect 1183 -295 1187 -291
rect 1232 -295 1236 -291
rect 77 -319 81 -315
rect 379 -318 383 -314
rect 559 -317 563 -313
rect 77 -327 81 -323
rect 379 -326 383 -322
rect 559 -325 563 -321
rect 559 -333 563 -329
rect 200 -341 204 -337
rect 559 -341 563 -337
rect 834 -348 838 -344
rect 77 -366 81 -362
rect 379 -359 383 -355
rect 834 -356 838 -352
rect 1253 -308 1257 -304
rect 77 -374 81 -370
rect 379 -367 383 -363
rect 763 -380 767 -376
rect 763 -388 767 -384
rect 914 -380 918 -376
rect -379 -393 -375 -389
rect -178 -394 -174 -390
rect 6 -398 10 -394
rect 6 -406 10 -402
rect 157 -398 161 -394
rect 914 -388 918 -384
rect 1145 -394 1149 -390
rect -348 -422 -344 -418
rect -299 -422 -295 -418
rect -389 -497 -385 -493
rect -340 -485 -336 -481
rect -291 -485 -287 -481
rect 157 -406 161 -402
rect 834 -412 838 -408
rect -147 -423 -143 -419
rect -98 -423 -94 -419
rect 834 -420 838 -416
rect 77 -430 81 -426
rect 77 -438 81 -434
rect 379 -430 383 -426
rect 379 -438 383 -434
rect 379 -446 383 -442
rect 555 -439 561 -433
rect -270 -498 -266 -494
rect -188 -498 -184 -494
rect -139 -486 -135 -482
rect -90 -486 -86 -482
rect 379 -454 383 -450
rect 77 -468 81 -464
rect 379 -462 383 -458
rect 77 -476 81 -472
rect -69 -499 -65 -495
rect 200 -490 204 -486
rect 379 -493 383 -489
rect 1176 -423 1180 -419
rect 1225 -423 1229 -419
rect 77 -516 81 -512
rect 379 -509 383 -505
rect 535 -501 539 -497
rect 1135 -498 1139 -494
rect 1184 -486 1188 -482
rect 1233 -486 1237 -482
rect 77 -524 81 -520
rect 379 -517 383 -513
rect 535 -509 539 -505
rect 6 -548 10 -544
rect 6 -556 10 -552
rect 157 -548 161 -544
rect 379 -547 383 -543
rect 1254 -499 1258 -495
rect 157 -556 161 -552
rect 379 -555 383 -551
rect 379 -563 383 -559
rect 535 -565 539 -561
rect -377 -583 -373 -579
rect 77 -580 81 -576
rect 535 -573 539 -569
rect -176 -584 -172 -580
rect 77 -588 81 -584
rect 535 -581 539 -577
rect 379 -596 383 -592
rect 535 -589 539 -585
rect 1147 -584 1151 -580
rect -346 -612 -342 -608
rect -297 -612 -293 -608
rect -387 -687 -383 -683
rect -338 -675 -334 -671
rect -289 -675 -285 -671
rect 379 -604 383 -600
rect 535 -597 539 -593
rect -145 -613 -141 -609
rect -96 -613 -92 -609
rect 77 -618 81 -614
rect 77 -626 81 -622
rect -268 -688 -264 -684
rect -186 -688 -182 -684
rect -137 -676 -133 -672
rect -88 -676 -84 -672
rect 200 -640 204 -636
rect 1178 -613 1182 -609
rect 1227 -613 1231 -609
rect -67 -689 -63 -685
rect 1137 -688 1141 -684
rect 1186 -676 1190 -672
rect 1235 -676 1239 -672
rect 1256 -689 1260 -685
<< metal1 >>
rect -397 192 -358 196
rect -391 166 -387 192
rect -353 195 -273 196
rect -353 192 -157 195
rect -379 183 -344 186
rect -383 166 -379 171
rect -348 158 -344 183
rect -338 158 -334 173
rect -348 154 -318 158
rect -357 145 -353 149
rect -357 141 -348 145
rect -352 139 -348 141
rect -340 101 -330 103
rect -340 99 -325 101
rect -393 75 -389 79
rect -375 72 -371 86
rect -363 87 -340 91
rect -363 72 -359 87
rect -329 84 -325 99
rect -322 91 -318 154
rect -310 139 -306 192
rect -277 191 -157 192
rect -310 135 -303 139
rect -277 133 -273 191
rect -190 165 -186 191
rect -152 191 -72 195
rect 383 191 422 195
rect -178 182 -143 185
rect -277 129 -253 133
rect -271 125 -267 129
rect -295 95 -280 99
rect -322 87 -291 91
rect -383 68 -359 72
rect -383 50 -379 68
rect -391 28 -387 30
rect -352 27 -348 44
rect -332 80 -325 84
rect -344 39 -340 44
rect -303 27 -299 44
rect -283 78 -280 95
rect -182 165 -178 170
rect -147 157 -143 182
rect -137 157 -133 172
rect -147 153 -117 157
rect -156 144 -152 148
rect -156 140 -147 144
rect -151 138 -147 140
rect -139 100 -129 102
rect -139 98 -124 100
rect -283 74 -270 78
rect -263 77 -259 85
rect -263 73 -229 77
rect -192 74 -188 78
rect -263 71 -259 73
rect -295 39 -291 44
rect -271 28 -267 51
rect -387 23 -271 27
rect -233 13 -229 73
rect -174 71 -170 85
rect -162 86 -139 90
rect -162 71 -158 86
rect -128 83 -124 98
rect -121 90 -117 153
rect -109 138 -105 191
rect -109 134 -102 138
rect -76 132 -72 191
rect 389 165 393 191
rect 427 191 507 195
rect 1127 191 1166 195
rect 401 182 436 185
rect -76 128 -52 132
rect -70 124 -66 128
rect -94 94 -79 98
rect -121 86 -90 90
rect -182 67 -158 71
rect -182 49 -178 67
rect -190 27 -186 29
rect -151 26 -147 43
rect -131 79 -124 83
rect -143 38 -139 43
rect -102 26 -98 43
rect -82 77 -79 94
rect -82 73 -69 77
rect -62 76 -58 84
rect 0 82 77 86
rect 85 82 89 93
rect 134 86 142 90
rect 196 86 285 90
rect -62 72 -46 76
rect -62 70 -58 72
rect -50 69 -46 72
rect 0 59 4 82
rect 85 78 94 82
rect 71 74 77 78
rect 138 74 142 86
rect -33 55 4 59
rect -94 38 -90 43
rect -70 26 -66 50
rect -186 22 -66 26
rect -33 13 -29 55
rect 0 54 4 55
rect 0 50 6 54
rect 14 50 18 61
rect 71 58 75 74
rect 134 70 156 74
rect 63 54 75 58
rect 125 54 137 58
rect 147 54 151 70
rect 14 46 23 50
rect -14 42 6 46
rect 67 42 75 54
rect 147 50 157 54
rect 165 50 169 62
rect 218 58 222 67
rect 285 58 289 86
rect 397 165 401 170
rect 432 157 436 182
rect 442 157 446 172
rect 432 153 462 157
rect 423 144 427 148
rect 423 140 432 144
rect 428 138 432 140
rect 440 100 450 102
rect 440 98 455 100
rect 387 74 391 78
rect 405 71 409 85
rect 417 86 440 90
rect 417 71 421 86
rect 451 83 455 98
rect 458 90 462 153
rect 470 138 474 191
rect 470 134 477 138
rect 503 132 507 191
rect 1133 165 1137 191
rect 1171 191 1251 195
rect 1145 182 1180 185
rect 503 128 527 132
rect 509 124 513 128
rect 485 94 500 98
rect 458 86 489 90
rect 214 54 222 58
rect 276 54 289 58
rect 165 46 174 50
rect 147 42 157 46
rect 218 42 222 54
rect -233 9 -29 13
rect 0 14 4 42
rect 63 38 85 42
rect 71 22 75 38
rect 71 18 77 22
rect 85 18 89 30
rect 134 22 142 26
rect 85 14 94 18
rect 0 10 77 14
rect -396 -1 -357 3
rect -390 -27 -386 -1
rect -352 2 -272 3
rect -352 -1 -156 2
rect -378 -10 -343 -7
rect -382 -27 -378 -22
rect -347 -35 -343 -10
rect -337 -35 -333 -20
rect -347 -39 -317 -35
rect -356 -48 -352 -44
rect -356 -52 -347 -48
rect -351 -54 -347 -52
rect -339 -92 -329 -90
rect -339 -94 -324 -92
rect -392 -118 -388 -114
rect -374 -121 -370 -107
rect -362 -106 -339 -102
rect -362 -121 -358 -106
rect -328 -109 -324 -94
rect -321 -102 -317 -39
rect -309 -54 -305 -1
rect -276 -2 -156 -1
rect -309 -58 -302 -54
rect -276 -60 -272 -2
rect -189 -28 -185 -2
rect -151 -2 -71 2
rect -177 -11 -142 -8
rect -276 -64 -252 -60
rect -270 -68 -266 -64
rect -294 -98 -279 -94
rect -321 -106 -290 -102
rect -382 -125 -358 -121
rect -382 -143 -378 -125
rect -390 -165 -386 -163
rect -351 -166 -347 -149
rect -331 -113 -324 -109
rect -343 -154 -339 -149
rect -302 -166 -298 -149
rect -282 -115 -279 -98
rect -181 -28 -177 -23
rect -146 -36 -142 -11
rect -136 -36 -132 -21
rect -146 -40 -116 -36
rect -155 -49 -151 -45
rect -155 -53 -146 -49
rect -150 -55 -146 -53
rect -138 -93 -128 -91
rect -138 -95 -123 -93
rect -282 -119 -269 -115
rect -262 -116 -258 -108
rect -262 -120 -225 -116
rect -191 -119 -187 -115
rect -262 -122 -258 -120
rect -294 -154 -290 -149
rect -270 -165 -266 -142
rect -270 -166 -269 -165
rect -386 -170 -269 -166
rect -229 -177 -225 -120
rect -173 -122 -169 -108
rect -161 -107 -138 -103
rect -161 -122 -157 -107
rect -127 -110 -123 -95
rect -120 -103 -116 -40
rect -108 -55 -104 -2
rect -108 -59 -101 -55
rect -75 -61 -71 -2
rect -33 -24 -29 9
rect 36 -16 40 10
rect 36 -20 77 -16
rect 85 -20 89 14
rect 138 10 142 22
rect 147 10 151 42
rect 214 38 236 42
rect 213 26 217 30
rect 285 26 289 54
rect 397 67 421 71
rect 397 49 401 67
rect 196 22 289 26
rect 389 26 393 29
rect 428 26 432 43
rect 448 79 455 83
rect 436 38 440 43
rect 477 26 481 43
rect 497 77 500 94
rect 1141 165 1145 170
rect 1176 157 1180 182
rect 1186 157 1190 172
rect 1176 153 1206 157
rect 1167 144 1171 148
rect 1167 140 1176 144
rect 1172 138 1176 140
rect 1184 100 1194 102
rect 1184 98 1199 100
rect 497 73 510 77
rect 517 76 521 84
rect 517 73 533 76
rect 1131 74 1135 78
rect 517 70 521 73
rect 1149 71 1153 85
rect 1161 86 1184 90
rect 1161 71 1165 86
rect 1195 83 1199 98
rect 1202 90 1206 153
rect 1214 138 1218 191
rect 1214 134 1221 138
rect 1247 132 1251 191
rect 1247 128 1271 132
rect 1253 124 1257 128
rect 1229 94 1244 98
rect 1202 86 1233 90
rect 1141 67 1165 71
rect 485 38 489 43
rect 509 26 513 50
rect 1141 49 1145 67
rect 1133 27 1137 29
rect 389 22 513 26
rect 1172 26 1176 43
rect 1192 79 1199 83
rect 1180 38 1184 43
rect 1221 26 1225 43
rect 1241 77 1244 94
rect 1241 73 1254 77
rect 1261 76 1265 84
rect 1261 72 1277 76
rect 1261 70 1265 72
rect 1229 38 1233 43
rect 1253 27 1257 50
rect 1137 22 1253 26
rect 134 6 156 10
rect 213 -12 217 22
rect 285 9 289 22
rect 431 9 435 22
rect 285 5 435 9
rect 1128 -2 1167 2
rect 134 -16 142 -12
rect 196 -16 217 -12
rect 85 -24 94 -20
rect -33 -28 77 -24
rect 85 -40 89 -24
rect 138 -28 142 -16
rect 757 -18 834 -14
rect 842 -18 846 -7
rect 891 -14 899 -10
rect 953 -14 1042 -10
rect 757 -23 761 -18
rect 842 -22 851 -18
rect 268 -27 761 -23
rect 134 -32 156 -28
rect 144 -38 148 -32
rect 268 -37 272 -27
rect 85 -43 94 -40
rect 144 -42 201 -38
rect 261 -41 275 -37
rect 85 -45 98 -43
rect 85 -47 221 -45
rect 85 -51 89 -47
rect 93 -49 221 -47
rect 295 -49 299 -45
rect -75 -65 -51 -61
rect -69 -69 -65 -65
rect 0 -67 77 -63
rect 85 -67 89 -56
rect 285 -58 289 -49
rect 134 -63 142 -59
rect 196 -63 285 -59
rect 320 -61 324 -27
rect 336 -31 340 -27
rect 373 -40 377 -27
rect 436 -40 444 -36
rect 498 -40 677 -36
rect 373 -44 379 -40
rect 387 -48 396 -44
rect 373 -52 379 -48
rect -93 -99 -78 -95
rect -120 -107 -89 -103
rect -181 -126 -157 -122
rect -181 -144 -177 -126
rect -189 -165 -185 -164
rect -150 -167 -146 -150
rect -130 -114 -123 -110
rect -142 -155 -138 -150
rect -101 -167 -97 -150
rect -81 -116 -78 -99
rect 0 -89 4 -67
rect 85 -71 94 -67
rect 71 -75 77 -71
rect 138 -75 142 -63
rect -81 -120 -68 -116
rect -61 -117 -57 -109
rect -20 -93 4 -89
rect -61 -121 -45 -117
rect -61 -123 -57 -121
rect -49 -124 -45 -121
rect -93 -155 -89 -150
rect -69 -167 -65 -143
rect -185 -170 -65 -167
rect -190 -171 -65 -170
rect -20 -173 -16 -93
rect 0 -95 4 -93
rect 0 -99 6 -95
rect 14 -99 18 -88
rect 71 -91 75 -75
rect 134 -79 156 -75
rect 63 -95 75 -91
rect 125 -95 137 -91
rect 147 -95 151 -79
rect 14 -103 23 -99
rect 0 -107 6 -103
rect 67 -107 75 -95
rect 147 -99 157 -95
rect 165 -99 169 -87
rect 218 -91 222 -82
rect 285 -91 289 -63
rect 373 -78 377 -52
rect 387 -61 391 -48
rect 440 -52 444 -40
rect 673 -43 677 -40
rect 603 -48 611 -44
rect 665 -48 673 -44
rect 757 -46 761 -27
rect 828 -26 834 -22
rect 895 -26 899 -14
rect 522 -52 546 -48
rect 436 -56 458 -52
rect 498 -56 526 -52
rect 554 -56 563 -52
rect 607 -54 611 -48
rect 757 -50 763 -46
rect 771 -50 775 -39
rect 828 -42 832 -26
rect 891 -30 913 -26
rect 820 -46 832 -42
rect 882 -46 894 -42
rect 904 -46 908 -30
rect 533 -60 546 -56
rect 533 -68 537 -60
rect 465 -72 537 -68
rect 555 -69 559 -56
rect 607 -59 616 -54
rect 771 -54 780 -50
rect 757 -58 763 -54
rect 824 -58 832 -46
rect 904 -50 914 -46
rect 922 -50 926 -38
rect 975 -42 979 -33
rect 1042 -42 1046 -14
rect 971 -46 979 -42
rect 1033 -46 1046 -42
rect 922 -54 931 -50
rect 904 -58 914 -54
rect 975 -58 979 -46
rect 607 -60 613 -59
rect 603 -64 613 -60
rect 618 -64 625 -60
rect 757 -78 761 -58
rect 820 -62 842 -58
rect 301 -82 761 -78
rect 828 -78 832 -62
rect 828 -82 834 -78
rect 842 -82 846 -70
rect 891 -78 899 -74
rect 757 -86 761 -82
rect 842 -86 851 -82
rect 683 -90 742 -86
rect 757 -90 834 -86
rect 214 -95 222 -91
rect 276 -95 289 -91
rect 165 -103 174 -99
rect 147 -107 157 -103
rect 218 -107 222 -95
rect 0 -124 4 -107
rect 63 -111 85 -107
rect 71 -127 75 -111
rect 0 -135 4 -129
rect 71 -131 77 -127
rect 85 -131 89 -119
rect 134 -127 142 -123
rect 85 -135 94 -131
rect 0 -139 77 -135
rect 36 -165 40 -139
rect 36 -169 77 -165
rect 85 -169 89 -135
rect 138 -139 142 -127
rect 147 -139 151 -107
rect 214 -111 236 -107
rect 213 -123 217 -119
rect 285 -123 289 -95
rect 196 -127 289 -123
rect 294 -95 460 -91
rect 134 -143 156 -139
rect 213 -161 217 -127
rect 294 -132 298 -95
rect 134 -165 142 -161
rect 196 -165 217 -161
rect 249 -136 298 -132
rect 85 -173 94 -169
rect -20 -177 77 -173
rect -229 -181 -16 -177
rect -398 -189 -359 -185
rect -392 -215 -388 -189
rect -354 -186 -274 -185
rect -354 -189 -158 -186
rect -380 -198 -345 -195
rect -384 -215 -380 -210
rect -349 -223 -345 -198
rect -339 -223 -335 -208
rect -349 -227 -319 -223
rect -358 -236 -354 -232
rect -358 -240 -349 -236
rect -353 -242 -349 -240
rect -341 -280 -331 -278
rect -341 -282 -326 -280
rect -394 -306 -390 -302
rect -376 -309 -372 -295
rect -364 -294 -341 -290
rect -364 -309 -360 -294
rect -330 -297 -326 -282
rect -323 -290 -319 -227
rect -311 -242 -307 -189
rect -278 -190 -158 -189
rect -311 -246 -304 -242
rect -278 -248 -274 -190
rect -191 -216 -187 -190
rect -153 -190 -73 -186
rect -179 -199 -144 -196
rect -278 -252 -254 -248
rect -272 -256 -268 -252
rect -296 -286 -281 -282
rect -323 -294 -292 -290
rect -384 -313 -360 -309
rect -384 -331 -380 -313
rect -392 -353 -388 -351
rect -353 -354 -349 -337
rect -333 -301 -326 -297
rect -345 -342 -341 -337
rect -304 -354 -300 -337
rect -284 -303 -281 -286
rect -183 -216 -179 -211
rect -148 -224 -144 -199
rect -138 -224 -134 -209
rect -148 -228 -118 -224
rect -157 -237 -153 -233
rect -157 -241 -148 -237
rect -152 -243 -148 -241
rect -140 -281 -130 -279
rect -140 -283 -125 -281
rect -284 -307 -271 -303
rect -264 -304 -260 -296
rect -264 -308 -247 -304
rect -193 -307 -189 -303
rect -264 -310 -260 -308
rect -296 -342 -292 -337
rect -272 -353 -268 -330
rect -272 -354 -271 -353
rect -388 -358 -271 -354
rect -251 -367 -247 -308
rect -175 -310 -171 -296
rect -163 -295 -140 -291
rect -163 -310 -159 -295
rect -129 -298 -125 -283
rect -122 -291 -118 -228
rect -110 -243 -106 -190
rect -110 -247 -103 -243
rect -77 -249 -73 -190
rect 85 -194 89 -173
rect 138 -177 142 -165
rect 249 -173 253 -136
rect 305 -143 310 -108
rect 389 -109 393 -106
rect 555 -109 559 -98
rect 320 -135 324 -109
rect 389 -113 582 -109
rect 320 -139 379 -135
rect 389 -139 393 -113
rect 441 -127 564 -123
rect 441 -131 445 -127
rect 437 -135 453 -131
rect 389 -143 397 -139
rect 305 -147 379 -143
rect 201 -177 253 -173
rect 268 -176 281 -172
rect 134 -181 156 -177
rect 144 -187 148 -181
rect 201 -187 205 -177
rect 268 -186 272 -176
rect 277 -177 281 -176
rect 144 -191 201 -187
rect 261 -190 275 -186
rect 85 -198 221 -194
rect 295 -198 299 -194
rect 0 -217 77 -213
rect 85 -217 89 -206
rect 285 -208 289 -198
rect 134 -213 142 -209
rect 196 -213 285 -209
rect 0 -237 4 -217
rect 85 -221 94 -217
rect 71 -225 77 -221
rect 138 -225 142 -213
rect -22 -241 4 -237
rect -77 -253 -53 -249
rect -71 -257 -67 -253
rect -95 -287 -80 -283
rect -122 -295 -91 -291
rect -183 -314 -159 -310
rect -183 -332 -179 -314
rect -191 -354 -187 -352
rect -152 -355 -148 -338
rect -132 -302 -125 -298
rect -144 -343 -140 -338
rect -103 -355 -99 -338
rect -83 -304 -80 -287
rect -83 -308 -70 -304
rect -63 -305 -59 -297
rect -63 -309 -47 -305
rect -63 -311 -59 -309
rect -51 -312 -47 -309
rect -22 -323 -18 -241
rect 0 -245 4 -241
rect 0 -249 6 -245
rect 14 -249 18 -238
rect 71 -241 75 -225
rect 134 -229 156 -225
rect 63 -245 75 -241
rect 125 -245 137 -241
rect 147 -245 151 -229
rect 14 -253 23 -249
rect 0 -257 6 -253
rect 67 -257 75 -245
rect 147 -249 157 -245
rect 165 -249 169 -237
rect 218 -241 222 -232
rect 285 -241 289 -213
rect 305 -217 310 -147
rect 332 -155 379 -151
rect 389 -155 393 -143
rect 441 -147 445 -135
rect 437 -151 445 -147
rect 560 -151 564 -127
rect 332 -228 336 -155
rect 389 -159 397 -155
rect 513 -159 519 -155
rect 560 -155 568 -151
rect 578 -155 582 -113
rect 738 -123 742 -90
rect 842 -101 846 -86
rect 895 -90 899 -78
rect 904 -90 908 -58
rect 971 -62 993 -58
rect 970 -74 974 -70
rect 1042 -74 1046 -46
rect 953 -78 1046 -74
rect 1134 -28 1138 -2
rect 1172 -2 1252 2
rect 1146 -11 1181 -8
rect 891 -94 913 -90
rect 970 -101 974 -78
rect 1142 -28 1146 -23
rect 1177 -36 1181 -11
rect 1187 -36 1191 -21
rect 1177 -40 1207 -36
rect 1168 -49 1172 -45
rect 1168 -53 1177 -49
rect 1173 -55 1177 -53
rect 1185 -93 1195 -91
rect 1185 -95 1200 -93
rect 738 -127 834 -123
rect 842 -127 846 -116
rect 891 -123 899 -119
rect 953 -123 1042 -119
rect 1132 -119 1136 -115
rect 1150 -122 1154 -108
rect 1162 -107 1185 -103
rect 1162 -122 1166 -107
rect 1196 -110 1200 -95
rect 1203 -103 1207 -40
rect 1215 -55 1219 -2
rect 1215 -59 1222 -55
rect 1248 -61 1252 -2
rect 1248 -65 1272 -61
rect 1254 -69 1258 -65
rect 1230 -99 1245 -95
rect 1203 -107 1234 -103
rect 630 -147 634 -139
rect 626 -151 642 -147
rect 578 -159 586 -155
rect 344 -184 349 -182
rect 344 -188 379 -184
rect 389 -188 393 -159
rect 519 -180 523 -159
rect 436 -184 444 -180
rect 498 -184 523 -180
rect 543 -163 568 -159
rect 387 -192 396 -188
rect 373 -196 379 -192
rect 373 -228 377 -196
rect 389 -206 393 -192
rect 440 -196 444 -184
rect 543 -196 547 -163
rect 436 -200 458 -196
rect 498 -200 547 -196
rect 560 -171 568 -167
rect 578 -171 582 -159
rect 630 -163 634 -151
rect 757 -155 761 -127
rect 842 -131 851 -127
rect 828 -135 834 -131
rect 895 -135 899 -123
rect 757 -159 763 -155
rect 771 -159 775 -148
rect 828 -151 832 -135
rect 891 -139 913 -135
rect 820 -155 832 -151
rect 882 -155 894 -151
rect 904 -155 908 -139
rect 771 -163 780 -159
rect 626 -167 634 -163
rect 757 -167 763 -163
rect 824 -167 832 -155
rect 904 -159 914 -155
rect 922 -159 926 -147
rect 975 -151 979 -142
rect 1042 -151 1046 -123
rect 1142 -126 1166 -122
rect 1142 -144 1146 -126
rect 971 -155 979 -151
rect 1033 -155 1046 -151
rect 922 -163 931 -159
rect 904 -167 914 -163
rect 975 -167 979 -155
rect 389 -210 418 -206
rect 560 -219 564 -171
rect 578 -175 586 -171
rect 630 -180 634 -167
rect 702 -175 712 -171
rect 757 -195 761 -167
rect 820 -171 842 -167
rect 828 -187 832 -171
rect 828 -191 834 -187
rect 842 -191 846 -179
rect 891 -187 899 -183
rect 842 -195 851 -191
rect 757 -196 834 -195
rect 399 -223 564 -219
rect 732 -199 834 -196
rect 732 -200 772 -199
rect 300 -232 588 -228
rect 732 -228 736 -200
rect 842 -210 846 -195
rect 895 -199 899 -187
rect 904 -199 908 -167
rect 971 -171 993 -167
rect 970 -183 974 -179
rect 1042 -183 1046 -155
rect 1134 -166 1138 -164
rect 1173 -167 1177 -150
rect 1193 -114 1200 -110
rect 1181 -155 1185 -150
rect 1222 -167 1226 -150
rect 1242 -116 1245 -99
rect 1242 -120 1255 -116
rect 1262 -117 1266 -109
rect 1262 -121 1278 -117
rect 1262 -123 1266 -121
rect 1230 -155 1234 -150
rect 1254 -166 1258 -143
rect 1254 -167 1255 -166
rect 1138 -171 1255 -167
rect 953 -187 1046 -183
rect 891 -203 913 -199
rect 970 -210 974 -187
rect 1126 -190 1165 -186
rect 1132 -216 1136 -190
rect 1170 -190 1250 -186
rect 1144 -199 1179 -196
rect 593 -232 736 -228
rect 214 -245 222 -241
rect 276 -245 289 -241
rect 165 -253 174 -249
rect 147 -257 157 -253
rect 218 -257 222 -245
rect 0 -285 4 -257
rect 63 -261 85 -257
rect 71 -277 75 -261
rect 71 -281 77 -277
rect 85 -281 89 -269
rect 134 -277 142 -273
rect 0 -289 15 -285
rect 85 -285 94 -281
rect 20 -289 77 -285
rect 45 -315 49 -289
rect 45 -319 77 -315
rect 85 -319 89 -285
rect 138 -289 142 -277
rect 147 -289 151 -257
rect 214 -261 236 -257
rect 213 -273 217 -269
rect 285 -273 289 -245
rect 196 -277 289 -273
rect 353 -268 357 -232
rect 363 -252 368 -250
rect 363 -256 379 -252
rect 386 -256 390 -244
rect 720 -243 725 -241
rect 757 -237 834 -233
rect 842 -237 846 -226
rect 891 -233 899 -229
rect 953 -233 1042 -229
rect 757 -243 761 -237
rect 842 -241 851 -237
rect 720 -247 761 -243
rect 436 -252 452 -248
rect 532 -252 557 -248
rect 386 -260 396 -256
rect 374 -264 379 -260
rect 353 -272 379 -268
rect 386 -272 390 -260
rect 440 -264 444 -252
rect 436 -268 444 -264
rect 134 -293 156 -289
rect 213 -311 217 -277
rect 134 -315 142 -311
rect 196 -315 217 -311
rect 256 -293 307 -289
rect 85 -323 94 -319
rect -22 -327 77 -323
rect -95 -343 -91 -338
rect -71 -355 -67 -331
rect -187 -359 -67 -355
rect -22 -367 -18 -327
rect 85 -341 89 -323
rect 138 -327 142 -315
rect 256 -323 260 -293
rect 319 -314 323 -283
rect 353 -306 357 -272
rect 386 -276 396 -272
rect 367 -280 379 -276
rect 367 -296 371 -280
rect 353 -310 379 -306
rect 389 -310 393 -276
rect 440 -280 444 -268
rect 436 -284 444 -280
rect 532 -284 536 -280
rect 441 -302 445 -294
rect 437 -306 453 -302
rect 513 -306 549 -302
rect 389 -314 397 -310
rect 319 -318 379 -314
rect 207 -327 260 -323
rect 267 -326 356 -322
rect 134 -331 156 -327
rect 207 -329 211 -327
rect 144 -337 148 -331
rect 200 -333 211 -329
rect 200 -337 204 -333
rect 267 -336 271 -326
rect 144 -341 200 -337
rect 260 -340 274 -336
rect 85 -342 94 -341
rect 85 -344 99 -342
rect 85 -346 220 -344
rect 85 -350 89 -346
rect 94 -348 220 -346
rect 294 -348 298 -344
rect -251 -371 -18 -367
rect 0 -366 77 -362
rect 85 -366 89 -355
rect 285 -357 289 -348
rect 134 -362 142 -358
rect 196 -362 285 -358
rect -397 -380 -358 -376
rect -391 -406 -387 -380
rect -353 -377 -273 -376
rect -353 -380 -157 -377
rect -379 -389 -344 -386
rect -383 -406 -379 -401
rect -348 -414 -344 -389
rect -338 -414 -334 -399
rect -348 -418 -318 -414
rect -357 -427 -353 -423
rect -357 -431 -348 -427
rect -352 -433 -348 -431
rect -340 -471 -330 -469
rect -340 -473 -325 -471
rect -393 -497 -389 -493
rect -375 -500 -371 -486
rect -363 -485 -340 -481
rect -363 -500 -359 -485
rect -329 -488 -325 -473
rect -322 -481 -318 -418
rect -310 -433 -306 -380
rect -277 -381 -157 -380
rect -310 -437 -303 -433
rect -277 -439 -273 -381
rect -190 -407 -186 -381
rect -152 -381 -72 -377
rect -178 -390 -143 -387
rect -277 -443 -253 -439
rect -271 -447 -267 -443
rect -295 -477 -280 -473
rect -322 -485 -291 -481
rect -383 -504 -359 -500
rect -383 -522 -379 -504
rect -391 -544 -387 -542
rect -352 -545 -348 -528
rect -332 -492 -325 -488
rect -344 -533 -340 -528
rect -303 -545 -299 -528
rect -283 -494 -280 -477
rect -182 -407 -178 -402
rect -147 -415 -143 -390
rect -137 -415 -133 -400
rect -147 -419 -117 -415
rect -156 -428 -152 -424
rect -156 -432 -147 -428
rect -151 -434 -147 -432
rect -139 -472 -129 -470
rect -139 -474 -124 -472
rect -283 -498 -270 -494
rect -263 -495 -259 -487
rect -263 -499 -237 -495
rect -192 -498 -188 -494
rect -263 -501 -259 -499
rect -295 -533 -291 -528
rect -271 -544 -267 -521
rect -271 -545 -269 -544
rect -387 -549 -269 -545
rect -241 -558 -237 -499
rect -174 -501 -170 -487
rect -162 -486 -139 -482
rect -162 -501 -158 -486
rect -128 -489 -124 -474
rect -121 -482 -117 -419
rect -109 -434 -105 -381
rect -109 -438 -102 -434
rect -76 -440 -72 -381
rect 0 -383 4 -366
rect 85 -370 94 -366
rect 71 -374 77 -370
rect 138 -374 142 -362
rect -21 -387 4 -383
rect -76 -444 -52 -440
rect -70 -448 -66 -444
rect -94 -478 -79 -474
rect -121 -486 -90 -482
rect -182 -505 -158 -501
rect -182 -523 -178 -505
rect -190 -545 -186 -543
rect -151 -546 -147 -529
rect -131 -493 -124 -489
rect -143 -534 -139 -529
rect -102 -546 -98 -529
rect -82 -495 -79 -478
rect -21 -472 -17 -387
rect 0 -394 4 -387
rect 0 -398 6 -394
rect 14 -398 18 -387
rect 71 -390 75 -374
rect 134 -378 156 -374
rect 63 -394 75 -390
rect 125 -394 137 -390
rect 147 -394 151 -378
rect 14 -402 23 -398
rect 0 -406 6 -402
rect 67 -406 75 -394
rect 147 -398 157 -394
rect 165 -398 169 -386
rect 218 -390 222 -381
rect 285 -390 289 -362
rect 214 -394 222 -390
rect 276 -394 289 -390
rect 165 -402 174 -398
rect 147 -406 157 -402
rect 218 -406 222 -394
rect 0 -434 4 -406
rect 63 -410 85 -406
rect 71 -426 75 -410
rect 71 -430 77 -426
rect 85 -430 89 -418
rect 134 -426 142 -422
rect 0 -438 11 -434
rect 85 -434 94 -430
rect 16 -438 77 -434
rect 45 -464 49 -438
rect 45 -468 77 -464
rect 85 -468 89 -434
rect 138 -438 142 -426
rect 147 -438 151 -406
rect 214 -410 236 -406
rect 213 -422 217 -418
rect 285 -422 289 -394
rect 196 -426 289 -422
rect 134 -442 156 -438
rect 213 -460 217 -426
rect 303 -448 307 -326
rect 352 -355 356 -326
rect 363 -326 379 -322
rect 389 -326 393 -314
rect 441 -318 445 -306
rect 437 -322 445 -318
rect 545 -321 549 -306
rect 553 -313 557 -252
rect 757 -265 761 -247
rect 828 -245 834 -241
rect 895 -245 899 -233
rect 757 -269 763 -265
rect 771 -269 775 -258
rect 828 -261 832 -245
rect 891 -249 913 -245
rect 820 -265 832 -261
rect 882 -265 894 -261
rect 904 -265 908 -249
rect 771 -273 780 -269
rect 588 -297 592 -276
rect 757 -277 763 -273
rect 824 -277 832 -265
rect 904 -269 914 -265
rect 922 -269 926 -257
rect 975 -261 979 -252
rect 1042 -261 1046 -233
rect 971 -265 979 -261
rect 1033 -265 1046 -261
rect 922 -273 931 -269
rect 904 -277 914 -273
rect 975 -277 979 -265
rect 601 -296 605 -278
rect 757 -301 761 -277
rect 820 -281 842 -277
rect 828 -297 832 -281
rect 828 -301 834 -297
rect 842 -301 846 -289
rect 891 -297 899 -293
rect 737 -305 761 -301
rect 842 -305 851 -301
rect 553 -317 559 -313
rect 566 -317 570 -305
rect 616 -313 632 -309
rect 566 -321 576 -317
rect 545 -325 559 -321
rect 363 -331 367 -326
rect 389 -330 397 -326
rect 513 -330 515 -326
rect 389 -341 393 -330
rect 546 -333 559 -329
rect 566 -333 570 -321
rect 620 -325 624 -313
rect 616 -329 624 -325
rect 566 -337 576 -333
rect 547 -339 559 -337
rect 389 -342 539 -341
rect 378 -345 539 -342
rect 552 -341 559 -339
rect 378 -346 393 -345
rect 352 -359 379 -355
rect 389 -359 393 -346
rect 535 -350 539 -345
rect 566 -350 570 -337
rect 620 -341 624 -329
rect 616 -345 624 -341
rect 712 -345 722 -341
rect 436 -355 444 -351
rect 498 -355 506 -351
rect 535 -354 570 -350
rect 620 -355 624 -345
rect 387 -363 396 -359
rect 372 -367 379 -363
rect 440 -367 444 -355
rect 372 -377 376 -367
rect 436 -371 458 -367
rect 498 -371 528 -367
rect 737 -377 741 -305
rect 757 -309 834 -305
rect 842 -320 846 -305
rect 895 -309 899 -297
rect 904 -309 908 -277
rect 971 -281 993 -277
rect 970 -293 974 -289
rect 1042 -293 1046 -265
rect 953 -297 1046 -293
rect 1140 -216 1144 -211
rect 1175 -224 1179 -199
rect 1185 -224 1189 -209
rect 1175 -228 1205 -224
rect 1166 -237 1170 -233
rect 1166 -241 1175 -237
rect 1171 -243 1175 -241
rect 1183 -281 1193 -279
rect 1183 -283 1198 -281
rect 891 -313 913 -309
rect 970 -320 974 -297
rect 1130 -307 1134 -303
rect 1148 -310 1152 -296
rect 1160 -295 1183 -291
rect 1160 -310 1164 -295
rect 1194 -298 1198 -283
rect 1201 -291 1205 -228
rect 1213 -243 1217 -190
rect 1213 -247 1220 -243
rect 1246 -249 1250 -190
rect 1246 -253 1270 -249
rect 1252 -257 1256 -253
rect 1228 -287 1243 -283
rect 1201 -295 1232 -291
rect 1140 -314 1164 -310
rect 1140 -332 1144 -314
rect 327 -381 741 -377
rect 757 -348 834 -344
rect 842 -348 846 -337
rect 891 -344 899 -340
rect 953 -344 1042 -340
rect 757 -355 761 -348
rect 842 -352 851 -348
rect 757 -360 758 -355
rect 828 -356 834 -352
rect 895 -356 899 -344
rect 757 -376 761 -360
rect 757 -380 763 -376
rect 771 -380 775 -369
rect 828 -372 832 -356
rect 891 -360 913 -356
rect 820 -376 832 -372
rect 882 -376 894 -372
rect 904 -376 908 -360
rect 771 -384 780 -380
rect 757 -388 763 -384
rect 824 -388 832 -376
rect 904 -380 914 -376
rect 922 -380 926 -368
rect 975 -372 979 -363
rect 1042 -372 1046 -344
rect 1132 -354 1136 -352
rect 1171 -355 1175 -338
rect 1191 -302 1198 -298
rect 1179 -343 1183 -338
rect 1220 -355 1224 -338
rect 1240 -304 1243 -287
rect 1240 -308 1253 -304
rect 1260 -305 1264 -297
rect 1260 -309 1276 -305
rect 1260 -311 1264 -309
rect 1228 -343 1232 -338
rect 1252 -354 1256 -331
rect 1252 -355 1253 -354
rect 1136 -359 1253 -355
rect 971 -376 979 -372
rect 1033 -376 1046 -372
rect 922 -384 931 -380
rect 904 -388 914 -384
rect 975 -388 979 -376
rect 340 -393 379 -389
rect 757 -397 761 -388
rect 820 -392 842 -388
rect 322 -401 761 -397
rect 134 -464 142 -460
rect 196 -464 217 -460
rect 85 -472 94 -468
rect -82 -499 -69 -495
rect -62 -496 -58 -488
rect -33 -476 77 -472
rect -62 -500 -46 -496
rect -62 -502 -58 -500
rect -50 -503 -46 -500
rect -94 -534 -90 -529
rect -70 -546 -66 -522
rect -186 -550 -66 -546
rect -33 -558 -29 -476
rect 85 -493 89 -472
rect 138 -476 142 -464
rect 207 -473 249 -469
rect 134 -480 156 -476
rect 144 -486 148 -480
rect 207 -482 211 -473
rect 200 -486 211 -482
rect 267 -475 291 -471
rect 267 -485 271 -475
rect 144 -490 200 -486
rect 260 -489 274 -485
rect 85 -497 220 -493
rect 294 -497 298 -493
rect 0 -516 77 -512
rect 85 -516 89 -505
rect 285 -507 289 -497
rect 134 -512 142 -508
rect 196 -512 285 -508
rect 0 -536 4 -516
rect 85 -520 94 -516
rect 71 -524 77 -520
rect 138 -524 142 -512
rect -241 -562 -29 -558
rect -24 -540 4 -536
rect -395 -570 -356 -566
rect -389 -596 -385 -570
rect -351 -567 -271 -566
rect -351 -570 -155 -567
rect -377 -579 -342 -576
rect -381 -596 -377 -591
rect -346 -604 -342 -579
rect -336 -604 -332 -589
rect -346 -608 -316 -604
rect -355 -617 -351 -613
rect -355 -621 -346 -617
rect -350 -623 -346 -621
rect -338 -661 -328 -659
rect -338 -663 -323 -661
rect -391 -687 -387 -683
rect -373 -690 -369 -676
rect -361 -675 -338 -671
rect -361 -690 -357 -675
rect -327 -678 -323 -663
rect -320 -671 -316 -608
rect -308 -623 -304 -570
rect -275 -571 -155 -570
rect -308 -627 -301 -623
rect -275 -629 -271 -571
rect -188 -597 -184 -571
rect -150 -571 -70 -567
rect -176 -580 -141 -577
rect -275 -633 -251 -629
rect -269 -637 -265 -633
rect -293 -667 -278 -663
rect -320 -675 -289 -671
rect -381 -694 -357 -690
rect -381 -712 -377 -694
rect -389 -734 -385 -732
rect -350 -735 -346 -718
rect -330 -682 -323 -678
rect -342 -723 -338 -718
rect -301 -735 -297 -718
rect -281 -684 -278 -667
rect -180 -597 -176 -592
rect -145 -605 -141 -580
rect -135 -605 -131 -590
rect -145 -609 -115 -605
rect -154 -618 -150 -614
rect -154 -622 -145 -618
rect -149 -624 -145 -622
rect -137 -662 -127 -660
rect -137 -664 -122 -662
rect -281 -688 -268 -684
rect -261 -685 -257 -677
rect -261 -689 -235 -685
rect -190 -688 -186 -684
rect -261 -691 -257 -689
rect -293 -723 -289 -718
rect -269 -734 -265 -711
rect -269 -735 -268 -734
rect -385 -739 -268 -735
rect -239 -750 -235 -689
rect -172 -691 -168 -677
rect -160 -676 -137 -672
rect -160 -691 -156 -676
rect -126 -679 -122 -664
rect -119 -672 -115 -609
rect -107 -624 -103 -571
rect -107 -628 -100 -624
rect -74 -630 -70 -571
rect -24 -622 -20 -540
rect 0 -544 4 -540
rect 0 -548 6 -544
rect 14 -548 18 -537
rect 71 -540 75 -524
rect 134 -528 156 -524
rect 63 -544 75 -540
rect 125 -544 137 -540
rect 147 -544 151 -528
rect 14 -552 23 -548
rect 0 -556 6 -552
rect 67 -556 75 -544
rect 147 -548 157 -544
rect 165 -548 169 -536
rect 218 -540 222 -531
rect 285 -540 289 -512
rect 214 -544 222 -540
rect 276 -544 289 -540
rect 165 -552 174 -548
rect 147 -556 157 -552
rect 218 -556 222 -544
rect 0 -584 4 -556
rect 63 -560 85 -556
rect 71 -576 75 -560
rect 71 -580 77 -576
rect 85 -580 89 -568
rect 134 -576 142 -572
rect 0 -588 15 -584
rect 85 -584 94 -580
rect 20 -588 77 -584
rect 32 -614 36 -588
rect 32 -618 77 -614
rect 85 -618 89 -584
rect 138 -588 142 -576
rect 147 -588 151 -556
rect 214 -560 236 -556
rect 213 -572 217 -568
rect 285 -572 289 -544
rect 196 -576 289 -572
rect 322 -526 326 -401
rect 345 -416 350 -414
rect 345 -420 360 -416
rect 356 -426 360 -420
rect 356 -430 379 -426
rect 388 -430 392 -412
rect 440 -414 580 -410
rect 440 -422 444 -414
rect 436 -426 452 -422
rect 337 -453 346 -449
rect 134 -592 156 -588
rect 213 -610 217 -576
rect 322 -592 326 -531
rect 334 -573 338 -475
rect 342 -551 346 -453
rect 356 -489 360 -430
rect 388 -434 396 -430
rect 375 -438 379 -434
rect 369 -446 379 -441
rect 388 -446 392 -434
rect 440 -438 444 -426
rect 557 -433 561 -432
rect 436 -442 444 -438
rect 561 -440 566 -436
rect 388 -450 396 -446
rect 377 -454 379 -450
rect 368 -462 379 -458
rect 388 -462 392 -450
rect 440 -454 444 -442
rect 561 -445 572 -440
rect 436 -458 444 -454
rect 388 -466 396 -462
rect 552 -466 558 -462
rect 388 -479 392 -466
rect 386 -483 392 -479
rect 441 -478 556 -474
rect 356 -493 379 -489
rect 386 -493 390 -483
rect 441 -485 445 -478
rect 436 -489 452 -485
rect 356 -543 360 -493
rect 386 -497 396 -493
rect 373 -509 379 -505
rect 386 -509 390 -497
rect 440 -501 444 -489
rect 541 -496 546 -488
rect 537 -497 546 -496
rect 539 -501 546 -497
rect 436 -505 444 -501
rect 386 -513 396 -509
rect 376 -517 379 -513
rect 356 -547 379 -543
rect 389 -547 393 -513
rect 440 -517 444 -505
rect 539 -509 541 -505
rect 536 -510 541 -509
rect 436 -521 444 -517
rect 532 -521 536 -517
rect 441 -539 445 -531
rect 437 -543 453 -539
rect 389 -551 397 -547
rect 342 -555 379 -551
rect 373 -563 379 -559
rect 389 -563 393 -551
rect 441 -555 445 -543
rect 437 -559 445 -555
rect 389 -564 397 -563
rect 388 -567 397 -564
rect 322 -596 379 -592
rect 388 -596 392 -567
rect 441 -577 445 -559
rect 517 -563 521 -521
rect 552 -537 556 -478
rect 567 -483 572 -445
rect 569 -488 572 -483
rect 576 -519 580 -414
rect 757 -416 761 -401
rect 828 -408 832 -392
rect 828 -412 834 -408
rect 842 -412 846 -400
rect 891 -408 899 -404
rect 842 -416 851 -412
rect 757 -420 834 -416
rect 842 -431 846 -416
rect 895 -420 899 -408
rect 904 -420 908 -388
rect 971 -392 993 -388
rect 970 -404 974 -400
rect 1042 -404 1046 -376
rect 1127 -381 1166 -377
rect 953 -408 1046 -404
rect 1133 -407 1137 -381
rect 1171 -381 1251 -377
rect 1145 -390 1180 -387
rect 891 -424 913 -420
rect 970 -431 974 -408
rect 1141 -407 1145 -402
rect 1176 -415 1180 -390
rect 1186 -415 1190 -400
rect 1176 -419 1206 -415
rect 1167 -428 1171 -424
rect 1167 -432 1176 -428
rect 1172 -434 1176 -432
rect 1184 -472 1194 -470
rect 1184 -474 1199 -472
rect 590 -496 631 -492
rect 1131 -498 1135 -494
rect 1149 -501 1153 -487
rect 1161 -486 1184 -482
rect 1161 -501 1165 -486
rect 1195 -489 1199 -474
rect 1202 -482 1206 -419
rect 1214 -434 1218 -381
rect 1214 -438 1221 -434
rect 1247 -440 1251 -381
rect 1247 -444 1271 -440
rect 1253 -448 1257 -444
rect 1229 -478 1244 -474
rect 1202 -486 1233 -482
rect 513 -567 521 -563
rect 526 -541 556 -537
rect 563 -523 580 -519
rect 1141 -505 1165 -501
rect 1141 -523 1145 -505
rect 526 -569 530 -541
rect 563 -548 567 -523
rect 1133 -545 1137 -543
rect 535 -552 567 -548
rect 596 -550 927 -546
rect 1172 -546 1176 -529
rect 1192 -493 1199 -489
rect 1180 -534 1184 -529
rect 1221 -546 1225 -529
rect 1241 -495 1244 -478
rect 1241 -499 1254 -495
rect 1261 -496 1265 -488
rect 1261 -500 1277 -496
rect 1261 -502 1265 -500
rect 1229 -534 1233 -529
rect 1253 -545 1257 -522
rect 1253 -546 1255 -545
rect 1137 -550 1255 -546
rect 535 -561 539 -552
rect 596 -557 600 -550
rect 592 -561 608 -557
rect 544 -569 552 -565
rect 526 -573 535 -569
rect 441 -581 535 -577
rect 544 -581 548 -569
rect 596 -573 600 -561
rect 592 -577 600 -573
rect 544 -585 552 -581
rect 436 -592 444 -588
rect 498 -592 505 -588
rect 517 -589 535 -585
rect 387 -600 396 -596
rect 360 -601 379 -600
rect 339 -604 379 -601
rect 339 -605 365 -604
rect 134 -614 142 -610
rect 196 -614 217 -610
rect 85 -622 94 -618
rect -24 -626 77 -622
rect -74 -634 -50 -630
rect -68 -638 -64 -634
rect -92 -668 -77 -664
rect -119 -676 -88 -672
rect -180 -695 -156 -691
rect -180 -713 -176 -695
rect -188 -735 -184 -733
rect -149 -736 -145 -719
rect -129 -683 -122 -679
rect -141 -724 -137 -719
rect -100 -736 -96 -719
rect -80 -685 -77 -668
rect -80 -689 -67 -685
rect -60 -686 -56 -678
rect -60 -690 -44 -686
rect -60 -692 -56 -690
rect -48 -693 -44 -690
rect -92 -724 -88 -719
rect -68 -736 -64 -712
rect -184 -740 -64 -736
rect -24 -750 -20 -626
rect 85 -643 89 -622
rect 138 -626 142 -614
rect 251 -616 301 -612
rect 134 -630 156 -626
rect 251 -627 255 -616
rect 297 -620 301 -616
rect 144 -636 148 -630
rect 200 -631 255 -627
rect 267 -625 280 -621
rect 200 -636 204 -631
rect 267 -635 271 -625
rect 388 -629 392 -600
rect 440 -604 444 -592
rect 517 -604 521 -589
rect 436 -608 458 -604
rect 498 -608 521 -604
rect 527 -597 535 -593
rect 544 -597 548 -585
rect 596 -589 600 -577
rect 592 -593 600 -589
rect 527 -621 531 -597
rect 460 -625 531 -621
rect 544 -601 552 -597
rect 708 -601 725 -597
rect 544 -629 548 -601
rect 388 -633 548 -629
rect 144 -640 200 -636
rect 260 -639 274 -635
rect 388 -636 392 -633
rect 382 -640 392 -636
rect 85 -647 220 -643
rect 294 -647 299 -643
rect 923 -684 927 -550
rect 1129 -571 1168 -567
rect 1135 -597 1139 -571
rect 1173 -571 1253 -567
rect 1147 -580 1182 -577
rect 1143 -597 1147 -592
rect 1178 -605 1182 -580
rect 1188 -605 1192 -590
rect 1178 -609 1208 -605
rect 1169 -618 1173 -614
rect 1169 -622 1178 -618
rect 1174 -624 1178 -622
rect 1186 -662 1196 -660
rect 1186 -664 1201 -662
rect 923 -688 1137 -684
rect 1151 -691 1155 -677
rect 1163 -676 1186 -672
rect 1163 -691 1167 -676
rect 1197 -679 1201 -664
rect 1204 -672 1208 -609
rect 1216 -624 1220 -571
rect 1216 -628 1223 -624
rect 1249 -630 1253 -571
rect 1249 -634 1273 -630
rect 1255 -638 1259 -634
rect 1231 -668 1246 -664
rect 1204 -676 1235 -672
rect 1143 -695 1167 -691
rect 1143 -713 1147 -695
rect 1135 -735 1139 -733
rect 1174 -736 1178 -719
rect 1194 -683 1201 -679
rect 1182 -724 1186 -719
rect 1223 -736 1227 -719
rect 1243 -685 1246 -668
rect 1243 -689 1256 -685
rect 1263 -686 1267 -678
rect 1263 -690 1279 -686
rect 1263 -692 1267 -690
rect 1231 -724 1235 -719
rect 1255 -735 1259 -712
rect 1255 -736 1256 -735
rect 1139 -740 1256 -736
rect -239 -754 -20 -750
<< m2contact >>
rect -402 192 -397 197
rect -358 191 -353 196
rect -338 173 -333 178
rect -358 149 -353 154
rect -330 101 -325 106
rect -398 75 -393 80
rect -299 154 -294 159
rect -157 190 -152 195
rect 378 191 383 196
rect -392 23 -387 28
rect -137 172 -132 177
rect -157 148 -152 153
rect -129 100 -124 105
rect -197 74 -192 79
rect -271 23 -266 28
rect -98 153 -93 158
rect 422 190 427 195
rect 1122 191 1127 196
rect -191 22 -186 27
rect 85 93 90 98
rect 285 86 290 91
rect -50 64 -45 69
rect 14 61 19 66
rect 137 54 142 59
rect 218 67 223 72
rect 164 62 169 67
rect -19 42 -14 47
rect 442 172 447 177
rect 422 148 427 153
rect 450 100 455 105
rect 382 74 387 79
rect 481 153 486 158
rect 1166 190 1171 195
rect 85 30 90 35
rect -401 -1 -396 4
rect -357 -2 -352 3
rect -337 -20 -332 -15
rect -357 -44 -352 -39
rect -329 -92 -324 -87
rect -397 -118 -392 -113
rect -298 -39 -293 -34
rect -156 -3 -151 2
rect -391 -170 -386 -165
rect -136 -21 -131 -16
rect -156 -45 -151 -40
rect -128 -93 -123 -88
rect -196 -119 -191 -114
rect -269 -170 -264 -165
rect -97 -40 -92 -35
rect 213 30 218 35
rect 1186 172 1191 177
rect 1166 148 1171 153
rect 1194 100 1199 105
rect 1126 74 1131 79
rect 1225 153 1230 158
rect 1132 22 1137 27
rect 1253 22 1258 27
rect 1123 -2 1128 3
rect 842 -7 847 -2
rect 1042 -14 1047 -9
rect 85 -56 90 -51
rect 285 -63 290 -58
rect 336 -36 341 -31
rect -190 -170 -185 -165
rect -49 -129 -44 -124
rect 14 -88 19 -83
rect 137 -95 142 -90
rect 218 -82 223 -77
rect 164 -87 169 -82
rect 320 -66 325 -61
rect 296 -82 301 -77
rect 673 -48 678 -43
rect 771 -39 776 -34
rect 894 -46 899 -41
rect 975 -33 980 -28
rect 921 -38 926 -33
rect 387 -66 392 -61
rect 460 -72 465 -67
rect 613 -64 618 -59
rect 555 -74 560 -69
rect 842 -70 847 -65
rect 678 -90 683 -85
rect 0 -129 5 -124
rect 85 -119 90 -114
rect 213 -119 218 -114
rect 460 -95 465 -90
rect 555 -98 560 -93
rect 305 -108 310 -103
rect -403 -189 -398 -184
rect -359 -190 -354 -185
rect -339 -208 -334 -203
rect -359 -232 -354 -227
rect -331 -280 -326 -275
rect -399 -306 -394 -301
rect -300 -227 -295 -222
rect -158 -191 -153 -186
rect -393 -358 -388 -353
rect -138 -209 -133 -204
rect -158 -233 -153 -228
rect -130 -281 -125 -276
rect -198 -307 -193 -302
rect -271 -358 -266 -353
rect -99 -228 -94 -223
rect 320 -109 325 -104
rect 387 -106 393 -101
rect 277 -182 282 -177
rect 85 -206 90 -201
rect 285 -213 290 -208
rect -192 -359 -187 -354
rect -51 -317 -46 -312
rect 14 -238 19 -233
rect 137 -245 142 -240
rect 218 -232 223 -227
rect 164 -237 169 -232
rect 305 -222 310 -217
rect 295 -232 300 -227
rect 519 -159 524 -154
rect 970 -70 975 -65
rect 1167 -3 1172 2
rect 1187 -21 1192 -16
rect 1167 -45 1172 -40
rect 1195 -93 1200 -88
rect 842 -116 847 -111
rect 1042 -123 1047 -118
rect 1127 -119 1132 -114
rect 1226 -40 1231 -35
rect 344 -182 349 -177
rect 771 -148 776 -143
rect 894 -155 899 -150
rect 975 -142 980 -137
rect 921 -147 926 -142
rect 418 -210 423 -205
rect 394 -223 399 -218
rect 712 -175 717 -170
rect 630 -185 635 -180
rect 842 -179 847 -174
rect 588 -232 593 -227
rect 970 -179 975 -174
rect 1133 -171 1138 -166
rect 1255 -171 1260 -166
rect 1121 -190 1126 -185
rect 1165 -191 1170 -186
rect 842 -226 847 -221
rect 85 -269 90 -264
rect 15 -289 20 -284
rect 213 -269 218 -264
rect 385 -244 390 -239
rect 363 -250 368 -245
rect 720 -241 725 -236
rect 1042 -233 1047 -228
rect 369 -264 374 -259
rect 319 -283 324 -278
rect 307 -293 312 -288
rect 367 -301 372 -296
rect 536 -284 541 -279
rect 85 -355 90 -350
rect 285 -362 290 -357
rect -402 -380 -397 -375
rect -358 -381 -353 -376
rect -338 -399 -333 -394
rect -358 -423 -353 -418
rect -330 -471 -325 -466
rect -398 -497 -393 -492
rect -299 -418 -294 -413
rect -157 -382 -152 -377
rect -392 -549 -387 -544
rect -137 -400 -132 -395
rect -157 -424 -152 -419
rect -129 -472 -124 -467
rect -197 -498 -192 -493
rect -269 -549 -264 -544
rect -98 -419 -93 -414
rect -191 -550 -186 -545
rect 14 -387 19 -382
rect 137 -394 142 -389
rect 218 -381 223 -376
rect 164 -386 169 -381
rect 85 -418 90 -413
rect 11 -438 16 -433
rect 213 -418 218 -413
rect 771 -258 776 -253
rect 894 -265 899 -260
rect 975 -252 980 -247
rect 921 -257 926 -252
rect 588 -276 593 -271
rect 601 -278 606 -273
rect 588 -302 593 -297
rect 601 -301 606 -296
rect 842 -289 847 -284
rect 363 -336 368 -331
rect 515 -333 520 -326
rect 541 -333 546 -328
rect 373 -346 378 -341
rect 547 -344 552 -339
rect 722 -345 727 -340
rect 506 -355 511 -350
rect 620 -360 625 -355
rect 322 -381 327 -376
rect 528 -371 533 -366
rect 970 -289 975 -284
rect 1185 -209 1190 -204
rect 1165 -233 1170 -228
rect 1193 -281 1198 -276
rect 1125 -307 1130 -302
rect 1224 -228 1229 -223
rect 842 -337 847 -332
rect 1042 -344 1047 -339
rect 758 -360 763 -355
rect 771 -369 776 -364
rect 894 -376 899 -371
rect 975 -363 980 -358
rect 921 -368 926 -363
rect 1131 -359 1136 -354
rect 1253 -359 1258 -354
rect 335 -393 340 -388
rect 379 -393 384 -388
rect 303 -453 308 -448
rect -50 -508 -45 -503
rect 249 -473 254 -468
rect 291 -475 296 -470
rect 85 -505 90 -500
rect 285 -512 290 -507
rect -400 -570 -395 -565
rect -356 -571 -351 -566
rect -336 -589 -331 -584
rect -356 -613 -351 -608
rect -328 -661 -323 -656
rect -396 -687 -391 -682
rect -297 -608 -292 -603
rect -155 -572 -150 -567
rect -390 -739 -385 -734
rect -135 -590 -130 -585
rect -155 -614 -150 -609
rect -127 -662 -122 -657
rect -195 -688 -190 -683
rect -268 -739 -263 -734
rect -96 -609 -91 -604
rect 14 -537 19 -532
rect 137 -544 142 -539
rect 218 -531 223 -526
rect 164 -536 169 -531
rect 85 -568 90 -563
rect 15 -588 20 -583
rect 213 -568 218 -563
rect 345 -414 350 -409
rect 387 -412 392 -407
rect 332 -453 337 -448
rect 334 -475 339 -470
rect 322 -531 327 -526
rect 364 -445 369 -440
rect 561 -436 566 -431
rect 372 -454 377 -449
rect 363 -462 368 -457
rect 558 -466 563 -461
rect 541 -488 546 -483
rect 371 -517 376 -512
rect 541 -510 546 -505
rect 536 -521 541 -516
rect 368 -563 373 -558
rect 334 -578 339 -573
rect 564 -488 569 -483
rect 842 -400 847 -395
rect 970 -400 975 -395
rect 1122 -381 1127 -376
rect 1166 -382 1171 -377
rect 1186 -400 1191 -395
rect 1166 -424 1171 -419
rect 1194 -472 1199 -467
rect 585 -496 590 -491
rect 631 -496 636 -491
rect 1126 -498 1131 -493
rect 1225 -419 1230 -414
rect 1132 -550 1137 -545
rect 1255 -550 1260 -545
rect 505 -592 510 -587
rect 334 -605 339 -600
rect -189 -740 -184 -735
rect -48 -698 -43 -693
rect 297 -625 302 -620
rect 455 -625 460 -620
rect 725 -601 730 -596
rect 377 -640 382 -635
rect 299 -647 304 -642
rect 1124 -571 1129 -566
rect 1168 -572 1173 -567
rect 1188 -590 1193 -585
rect 1168 -614 1173 -609
rect 1196 -662 1201 -657
rect 1227 -609 1232 -604
rect 1134 -740 1139 -735
rect 1256 -740 1261 -735
<< metal2 >>
rect -450 206 453 207
rect -450 203 1321 206
rect -450 17 -446 203
rect -426 192 -402 196
rect -357 154 -353 191
rect -338 178 -334 203
rect -330 154 -299 158
rect -330 106 -326 154
rect -156 153 -152 190
rect -137 177 -133 203
rect 442 202 1321 203
rect 373 191 378 195
rect -129 153 -98 157
rect -129 105 -125 153
rect 373 114 377 191
rect 423 153 427 190
rect 442 177 446 202
rect 1098 191 1122 195
rect 450 153 481 157
rect 1167 153 1171 190
rect 1186 177 1190 202
rect 64 110 377 114
rect 64 97 68 110
rect 450 105 454 153
rect 1194 153 1225 157
rect 1194 105 1198 153
rect 19 93 85 97
rect 90 93 98 97
rect -405 75 -398 79
rect -204 74 -197 78
rect -45 64 -38 68
rect -42 46 -38 64
rect 14 66 18 93
rect 94 67 98 93
rect 290 86 296 90
rect 356 74 382 78
rect 1079 74 1126 78
rect 356 71 360 74
rect 223 67 360 71
rect 94 63 164 67
rect -42 42 -19 46
rect 94 34 98 63
rect 90 30 98 34
rect 137 34 141 54
rect 137 30 213 34
rect -401 24 -392 28
rect -266 23 -191 27
rect -450 13 -132 17
rect -450 -174 -446 13
rect -426 -1 -401 3
rect -356 -39 -352 -2
rect -337 -15 -333 13
rect -329 -39 -298 -35
rect -329 -87 -325 -39
rect -155 -40 -151 -3
rect -136 -16 -132 13
rect 776 -7 842 -3
rect 847 -7 855 -3
rect -128 -40 -97 -36
rect 771 -34 775 -7
rect 851 -33 855 -7
rect 1047 -14 1053 -10
rect 1079 -29 1083 74
rect 1118 23 1132 27
rect 1317 16 1321 202
rect 1187 12 1321 16
rect 1098 -2 1123 2
rect 980 -33 1083 -29
rect -128 -88 -124 -40
rect 336 -42 340 -36
rect 851 -37 921 -33
rect 678 -48 683 -44
rect 19 -56 85 -52
rect 90 -56 98 -52
rect 14 -83 18 -56
rect 94 -82 98 -56
rect 290 -63 296 -59
rect 223 -82 296 -78
rect 94 -86 164 -82
rect -404 -118 -397 -114
rect -203 -119 -196 -115
rect 94 -115 98 -86
rect 296 -87 310 -82
rect 90 -119 98 -115
rect 137 -115 141 -95
rect 305 -103 310 -87
rect 320 -104 324 -66
rect 387 -101 391 -66
rect 613 -69 617 -64
rect 460 -90 464 -72
rect 613 -73 682 -69
rect 851 -66 855 -37
rect 1168 -40 1172 -3
rect 1187 -16 1191 12
rect 847 -70 855 -66
rect 1195 -40 1226 -36
rect 894 -66 898 -46
rect 894 -70 970 -66
rect 555 -93 559 -74
rect 678 -85 682 -73
rect 1195 -88 1199 -40
rect 137 -119 213 -115
rect 776 -116 842 -112
rect 847 -116 855 -112
rect -44 -129 0 -125
rect 525 -137 677 -133
rect 525 -150 529 -137
rect 771 -143 775 -116
rect 851 -142 855 -116
rect 1047 -123 1053 -119
rect 1119 -119 1127 -115
rect 980 -142 1057 -138
rect 851 -146 921 -142
rect 524 -159 529 -150
rect -401 -169 -391 -165
rect -264 -170 -190 -166
rect 319 -169 502 -165
rect -450 -178 -134 -174
rect -450 -363 -446 -178
rect -426 -189 -403 -185
rect -358 -227 -354 -190
rect -339 -203 -335 -178
rect -331 -227 -300 -223
rect -331 -275 -327 -227
rect -157 -228 -153 -191
rect -138 -204 -134 -178
rect 319 -178 323 -169
rect 498 -173 502 -169
rect 498 -177 533 -173
rect 717 -175 721 -171
rect 282 -182 344 -178
rect 19 -206 85 -202
rect 90 -206 98 -202
rect -130 -228 -99 -224
rect -130 -276 -126 -228
rect 14 -233 18 -206
rect 94 -232 98 -206
rect 290 -213 296 -209
rect 223 -232 295 -228
rect 94 -236 164 -232
rect 94 -265 98 -236
rect 305 -237 310 -222
rect 90 -269 98 -265
rect 137 -265 141 -245
rect 137 -269 213 -265
rect 319 -278 323 -182
rect 529 -189 533 -177
rect 851 -175 855 -146
rect 1053 -147 1057 -142
rect 1119 -147 1123 -119
rect 847 -179 855 -175
rect 1053 -151 1123 -147
rect 894 -175 898 -155
rect 1118 -166 1119 -165
rect 1118 -170 1133 -166
rect 894 -179 970 -175
rect 1317 -175 1321 12
rect 1185 -179 1321 -175
rect 635 -185 724 -181
rect 529 -193 605 -189
rect 347 -223 394 -219
rect 347 -288 352 -223
rect 363 -245 370 -241
rect 368 -246 370 -245
rect 418 -240 422 -210
rect 390 -244 422 -240
rect 363 -264 369 -259
rect 588 -271 592 -232
rect 601 -273 605 -193
rect 720 -236 724 -185
rect 1098 -190 1121 -186
rect 776 -226 842 -222
rect 847 -226 855 -222
rect 771 -253 775 -226
rect 851 -252 855 -226
rect 1166 -228 1170 -191
rect 1185 -204 1189 -179
rect 1047 -233 1053 -229
rect 1193 -228 1224 -224
rect 980 -252 1057 -248
rect 851 -256 921 -252
rect -406 -306 -399 -302
rect -205 -307 -198 -303
rect 15 -313 19 -289
rect 312 -293 352 -288
rect 536 -286 541 -284
rect 536 -290 722 -286
rect 851 -285 855 -256
rect 847 -289 855 -285
rect 894 -285 898 -265
rect 894 -289 970 -285
rect 536 -293 540 -290
rect -46 -317 19 -313
rect 332 -301 367 -297
rect 520 -297 540 -293
rect 332 -332 336 -301
rect 318 -336 363 -332
rect 520 -330 524 -297
rect 528 -333 541 -329
rect -401 -357 -393 -353
rect -266 -358 -192 -354
rect 19 -355 85 -351
rect 90 -355 98 -351
rect -450 -367 -133 -363
rect -450 -555 -446 -367
rect -426 -380 -402 -376
rect -357 -418 -353 -381
rect -338 -394 -334 -367
rect -330 -418 -299 -414
rect -330 -466 -326 -418
rect -156 -419 -152 -382
rect -137 -395 -133 -367
rect 14 -382 18 -355
rect 94 -381 98 -355
rect 290 -362 296 -358
rect 318 -377 322 -336
rect 223 -381 322 -377
rect 94 -385 164 -381
rect -129 -419 -98 -415
rect 94 -414 98 -385
rect 90 -418 98 -414
rect 293 -393 335 -389
rect 137 -414 141 -394
rect 137 -418 213 -414
rect -129 -467 -125 -419
rect 11 -443 15 -438
rect -6 -447 15 -443
rect -405 -497 -398 -493
rect -204 -498 -197 -494
rect -6 -504 -2 -447
rect 293 -451 297 -393
rect 345 -409 349 -336
rect 362 -346 373 -342
rect 362 -408 366 -346
rect 515 -351 519 -333
rect 511 -355 519 -351
rect 528 -366 532 -333
rect 547 -389 551 -344
rect 384 -393 551 -389
rect 362 -412 387 -408
rect 332 -440 336 -429
rect 588 -432 592 -302
rect 601 -419 605 -301
rect 722 -340 726 -290
rect 1053 -303 1057 -252
rect 1193 -276 1197 -228
rect 1053 -307 1125 -303
rect 776 -337 842 -333
rect 847 -337 855 -333
rect 625 -360 758 -356
rect 771 -364 775 -337
rect 851 -363 855 -337
rect 1047 -344 1053 -340
rect 1118 -354 1119 -353
rect 1118 -358 1131 -354
rect 980 -363 1057 -359
rect 851 -367 921 -363
rect 851 -396 855 -367
rect 847 -400 855 -396
rect 894 -396 898 -376
rect 894 -400 970 -396
rect 601 -423 635 -419
rect 566 -436 592 -432
rect 332 -444 364 -440
rect 249 -455 297 -451
rect 308 -453 332 -449
rect 347 -453 372 -449
rect 347 -454 358 -453
rect 249 -468 253 -455
rect 347 -460 352 -454
rect 319 -465 352 -460
rect 362 -462 363 -457
rect 296 -475 334 -471
rect -45 -508 -2 -504
rect 19 -505 85 -501
rect 90 -505 98 -501
rect 14 -532 18 -505
rect 94 -531 98 -505
rect 290 -512 296 -508
rect 362 -513 366 -462
rect 563 -466 598 -462
rect 546 -488 564 -483
rect 565 -496 585 -492
rect 565 -506 569 -496
rect 546 -510 569 -506
rect 594 -503 598 -466
rect 631 -491 635 -423
rect 1053 -494 1057 -363
rect 1317 -364 1321 -179
rect 1186 -368 1321 -364
rect 1098 -381 1122 -377
rect 1167 -419 1171 -382
rect 1186 -395 1190 -368
rect 1194 -419 1225 -415
rect 1194 -467 1198 -419
rect 1053 -498 1126 -494
rect 594 -507 728 -503
rect 362 -517 371 -513
rect 223 -531 322 -527
rect 94 -535 164 -531
rect -401 -548 -392 -544
rect -264 -549 -191 -545
rect -450 -559 -131 -555
rect -426 -570 -400 -566
rect -355 -608 -351 -571
rect -336 -584 -332 -559
rect -328 -608 -297 -604
rect -328 -656 -324 -608
rect -154 -609 -150 -572
rect -135 -585 -131 -559
rect 94 -564 98 -535
rect 90 -568 98 -564
rect 137 -564 141 -544
rect 303 -559 307 -531
rect 362 -557 366 -517
rect 594 -517 598 -507
rect 541 -521 598 -517
rect 1118 -545 1119 -544
rect 1118 -549 1132 -545
rect 1317 -556 1321 -368
rect 362 -558 369 -557
rect 362 -559 368 -558
rect 303 -563 368 -559
rect 1188 -560 1321 -556
rect 137 -568 213 -564
rect 1098 -571 1124 -567
rect -127 -609 -96 -605
rect -127 -657 -123 -609
rect -403 -687 -396 -683
rect -202 -688 -195 -684
rect 15 -694 19 -588
rect 334 -600 338 -578
rect 505 -614 509 -592
rect 730 -601 734 -597
rect 1169 -609 1173 -572
rect 1188 -585 1192 -560
rect 505 -618 572 -614
rect 1196 -609 1227 -605
rect 302 -625 455 -621
rect 364 -640 377 -636
rect 304 -648 308 -643
rect 1196 -657 1200 -609
rect -43 -698 19 -694
rect -401 -738 -390 -734
rect -263 -739 -189 -735
rect 1118 -735 1119 -734
rect 1118 -739 1134 -735
<< m3contact >>
rect -431 192 -426 197
rect 1093 191 1098 196
rect 14 93 19 98
rect 296 86 301 91
rect -406 23 -401 28
rect -431 -1 -426 4
rect 771 -7 776 -2
rect 1053 -14 1058 -9
rect 1113 22 1118 27
rect 1093 -2 1098 3
rect 336 -47 341 -42
rect 683 -48 688 -43
rect 14 -56 19 -51
rect 296 -63 301 -58
rect 771 -116 776 -111
rect 677 -137 682 -132
rect 1053 -123 1058 -118
rect -406 -170 -401 -165
rect -431 -189 -426 -184
rect 721 -175 726 -170
rect 14 -206 19 -201
rect 296 -213 301 -208
rect 305 -242 310 -237
rect 1113 -170 1118 -165
rect 370 -246 375 -241
rect 358 -264 363 -259
rect 1093 -190 1098 -185
rect 771 -226 776 -221
rect 1053 -233 1058 -228
rect 722 -290 727 -285
rect -406 -358 -401 -353
rect 14 -355 19 -350
rect -431 -380 -426 -375
rect 296 -362 301 -357
rect 332 -429 337 -424
rect 771 -337 776 -332
rect 1053 -344 1058 -339
rect 1113 -358 1118 -353
rect 314 -465 319 -460
rect 14 -505 19 -500
rect 296 -512 301 -507
rect 1093 -381 1098 -376
rect 728 -507 733 -502
rect -406 -549 -401 -544
rect -431 -570 -426 -565
rect 1113 -549 1118 -544
rect 1093 -571 1098 -566
rect 734 -601 739 -596
rect 572 -618 577 -613
rect 359 -640 364 -635
rect 304 -653 309 -648
rect -406 -739 -401 -734
rect 1113 -739 1118 -734
<< metal3 >>
rect -431 216 -6 220
rect -431 198 -427 216
rect -432 197 -425 198
rect -432 192 -431 197
rect -426 192 -425 197
rect -432 191 -425 192
rect -431 5 -427 191
rect -10 97 -6 216
rect 1092 196 1099 197
rect 1092 191 1093 196
rect 1098 191 1099 196
rect 1092 190 1099 191
rect 13 98 20 99
rect 13 97 14 98
rect -10 93 14 97
rect 19 93 20 98
rect -407 28 -400 29
rect -407 27 -406 28
rect -413 23 -406 27
rect -401 23 -400 28
rect -407 22 -400 23
rect -432 4 -425 5
rect -432 -1 -431 4
rect -426 -1 -425 4
rect -432 -2 -425 -1
rect -431 -183 -427 -2
rect -10 -52 -6 93
rect 13 92 20 93
rect 295 91 302 92
rect 295 86 296 91
rect 301 90 302 91
rect 301 86 312 90
rect 295 85 302 86
rect 1093 35 1097 190
rect 747 31 1097 35
rect 747 -3 751 31
rect 1093 4 1097 31
rect 1112 27 1119 28
rect 1112 26 1113 27
rect 1106 22 1113 26
rect 1118 22 1119 27
rect 1112 21 1119 22
rect 1092 3 1099 4
rect 770 -2 777 -1
rect 770 -3 771 -2
rect 747 -7 771 -3
rect 776 -7 777 -2
rect 1092 -2 1093 3
rect 1098 -2 1099 3
rect 1092 -3 1099 -2
rect 335 -42 342 -41
rect 335 -47 336 -42
rect 341 -47 342 -42
rect 335 -48 342 -47
rect 13 -51 20 -50
rect 13 -52 14 -51
rect -10 -56 14 -52
rect 19 -56 20 -51
rect 336 -51 342 -48
rect 682 -43 689 -42
rect 682 -48 683 -43
rect 688 -47 738 -43
rect 688 -48 689 -47
rect 682 -49 689 -48
rect -407 -165 -400 -164
rect -407 -166 -406 -165
rect -413 -170 -406 -166
rect -401 -170 -400 -165
rect -407 -171 -400 -170
rect -432 -184 -425 -183
rect -432 -189 -431 -184
rect -426 -189 -425 -184
rect -432 -190 -425 -189
rect -431 -374 -427 -190
rect -10 -202 -6 -56
rect 13 -57 20 -56
rect 295 -58 302 -57
rect 295 -63 296 -58
rect 301 -59 302 -58
rect 301 -63 312 -59
rect 295 -64 302 -63
rect 676 -132 683 -131
rect 734 -132 738 -47
rect 676 -137 677 -132
rect 682 -136 738 -132
rect 682 -137 683 -136
rect 676 -138 683 -137
rect 720 -170 727 -169
rect 734 -170 738 -136
rect 720 -175 721 -170
rect 726 -174 738 -170
rect 726 -175 727 -174
rect 720 -176 727 -175
rect 13 -201 20 -200
rect 13 -202 14 -201
rect -10 -206 14 -202
rect 19 -206 20 -201
rect -10 -351 -6 -206
rect 13 -207 20 -206
rect 295 -208 302 -207
rect 295 -213 296 -208
rect 301 -209 302 -208
rect 301 -213 312 -209
rect 295 -214 302 -213
rect 304 -237 311 -236
rect 304 -242 305 -237
rect 310 -242 311 -237
rect 304 -243 311 -242
rect 369 -241 376 -240
rect 305 -257 310 -243
rect 369 -246 370 -241
rect 375 -246 376 -241
rect 369 -247 376 -246
rect 305 -258 363 -257
rect 305 -259 364 -258
rect 305 -262 358 -259
rect 314 -327 319 -262
rect 357 -264 358 -262
rect 363 -264 364 -259
rect 357 -265 364 -264
rect 721 -285 728 -284
rect 734 -285 738 -174
rect 721 -290 722 -285
rect 727 -289 738 -285
rect 727 -290 728 -289
rect 721 -291 728 -290
rect 314 -332 328 -327
rect 13 -350 20 -349
rect 13 -351 14 -350
rect -407 -353 -400 -352
rect -407 -354 -406 -353
rect -413 -358 -406 -354
rect -401 -358 -400 -353
rect -407 -359 -400 -358
rect -10 -355 14 -351
rect 19 -355 20 -350
rect -432 -375 -425 -374
rect -432 -380 -431 -375
rect -426 -380 -425 -375
rect -432 -381 -425 -380
rect -431 -564 -427 -381
rect -10 -501 -6 -355
rect 13 -356 20 -355
rect 295 -357 302 -356
rect 295 -362 296 -357
rect 301 -358 302 -357
rect 301 -362 312 -358
rect 295 -363 302 -362
rect 323 -368 328 -332
rect 314 -373 328 -368
rect 314 -459 319 -373
rect 332 -423 337 -419
rect 331 -424 338 -423
rect 331 -429 332 -424
rect 337 -429 338 -424
rect 331 -430 338 -429
rect 313 -460 320 -459
rect 313 -465 314 -460
rect 319 -465 320 -460
rect 313 -466 320 -465
rect 13 -500 20 -499
rect 13 -501 14 -500
rect -10 -505 14 -501
rect 19 -505 20 -500
rect 734 -501 738 -289
rect -407 -544 -400 -543
rect -407 -545 -406 -544
rect -413 -549 -406 -545
rect -401 -549 -400 -544
rect -407 -550 -400 -549
rect -432 -565 -425 -564
rect -432 -570 -431 -565
rect -426 -570 -425 -565
rect -432 -571 -425 -570
rect -10 -679 -6 -505
rect 13 -506 20 -505
rect 727 -502 738 -501
rect 295 -507 302 -506
rect 727 -507 728 -502
rect 733 -507 738 -502
rect 295 -512 296 -507
rect 301 -508 302 -507
rect 301 -512 312 -508
rect 727 -508 738 -507
rect 295 -513 302 -512
rect 734 -595 738 -508
rect 747 -112 751 -7
rect 770 -8 777 -7
rect 1052 -9 1059 -8
rect 1052 -14 1053 -9
rect 1058 -10 1059 -9
rect 1058 -14 1069 -10
rect 1052 -15 1059 -14
rect 770 -111 777 -110
rect 770 -112 771 -111
rect 747 -116 771 -112
rect 776 -116 777 -111
rect 747 -222 751 -116
rect 770 -117 777 -116
rect 1052 -118 1059 -117
rect 1052 -123 1053 -118
rect 1058 -119 1059 -118
rect 1058 -123 1069 -119
rect 1052 -124 1059 -123
rect 1093 -184 1097 -3
rect 1112 -165 1119 -164
rect 1112 -166 1113 -165
rect 1106 -170 1113 -166
rect 1118 -170 1119 -165
rect 1112 -171 1119 -170
rect 1092 -185 1099 -184
rect 1092 -190 1093 -185
rect 1098 -190 1099 -185
rect 1092 -191 1099 -190
rect 770 -221 777 -220
rect 770 -222 771 -221
rect 747 -226 771 -222
rect 776 -226 777 -221
rect 747 -333 751 -226
rect 770 -227 777 -226
rect 1052 -228 1059 -227
rect 1052 -233 1053 -228
rect 1058 -229 1059 -228
rect 1058 -233 1069 -229
rect 1052 -234 1059 -233
rect 770 -332 777 -331
rect 770 -333 771 -332
rect 747 -337 771 -333
rect 776 -337 777 -332
rect 733 -596 740 -595
rect 733 -601 734 -596
rect 739 -601 740 -596
rect 733 -602 740 -601
rect 571 -613 578 -612
rect 734 -613 738 -602
rect 571 -618 572 -613
rect 577 -617 738 -613
rect 747 -616 751 -337
rect 770 -338 777 -337
rect 1052 -339 1059 -338
rect 1052 -344 1053 -339
rect 1058 -340 1059 -339
rect 1058 -344 1069 -340
rect 1052 -345 1059 -344
rect 1093 -375 1097 -191
rect 1112 -353 1119 -352
rect 1112 -354 1113 -353
rect 1106 -358 1113 -354
rect 1118 -358 1119 -353
rect 1112 -359 1119 -358
rect 1092 -376 1099 -375
rect 1092 -381 1093 -376
rect 1098 -381 1099 -376
rect 1092 -382 1099 -381
rect 1093 -565 1097 -382
rect 1112 -544 1119 -543
rect 1112 -545 1113 -544
rect 1106 -549 1113 -545
rect 1118 -549 1119 -544
rect 1112 -550 1119 -549
rect 1092 -566 1099 -565
rect 1092 -571 1093 -566
rect 1098 -571 1099 -566
rect 1092 -572 1099 -571
rect 747 -617 752 -616
rect 577 -618 578 -617
rect 571 -619 578 -618
rect 356 -635 365 -634
rect 352 -640 359 -635
rect 364 -640 365 -635
rect 352 -642 365 -640
rect 303 -648 309 -647
rect 303 -653 304 -648
rect 303 -654 309 -653
rect 304 -656 309 -654
rect 352 -679 356 -642
rect 734 -657 738 -617
rect 653 -661 738 -657
rect 748 -679 752 -617
rect -10 -683 752 -679
rect -407 -734 -400 -733
rect -407 -735 -406 -734
rect -413 -739 -406 -735
rect -401 -739 -400 -734
rect 1112 -734 1119 -733
rect 1112 -735 1113 -734
rect -407 -740 -400 -739
rect 1106 -739 1113 -735
rect 1118 -739 1119 -734
rect 1112 -740 1119 -739
<< m4contact >>
rect -418 22 -413 27
rect 312 86 317 91
rect 1101 21 1106 26
rect 336 -56 341 -51
rect -418 -171 -413 -166
rect 312 -63 317 -58
rect 312 -213 317 -208
rect 370 -240 375 -235
rect -418 -359 -413 -354
rect 312 -362 317 -357
rect 332 -419 337 -414
rect -418 -550 -413 -545
rect 312 -512 317 -507
rect 1069 -14 1074 -9
rect 1069 -123 1074 -118
rect 1101 -171 1106 -166
rect 1069 -233 1074 -228
rect 1069 -344 1074 -339
rect 1101 -359 1106 -354
rect 1101 -550 1106 -545
rect 304 -661 309 -656
rect 648 -661 653 -656
rect -418 -740 -413 -735
rect 1101 -740 1106 -735
<< metal4 >>
rect 312 91 316 92
rect -436 27 -432 28
rect -436 23 -418 27
rect -436 -166 -432 23
rect 312 -58 316 86
rect 1069 22 1101 26
rect 1069 -9 1073 22
rect 336 -59 341 -56
rect -436 -170 -418 -166
rect -436 -354 -432 -170
rect 312 -208 316 -63
rect 1069 -118 1073 -14
rect 1069 -166 1073 -123
rect 1069 -170 1101 -166
rect -436 -358 -418 -354
rect -436 -545 -432 -358
rect 312 -357 316 -213
rect 1069 -228 1073 -170
rect 365 -240 370 -236
rect 1069 -339 1073 -233
rect 1069 -354 1073 -344
rect 1069 -358 1101 -354
rect 312 -507 316 -362
rect 332 -414 336 -410
rect -436 -549 -418 -545
rect -436 -735 -432 -549
rect 312 -656 316 -512
rect 1069 -545 1073 -358
rect 1069 -549 1101 -545
rect 309 -657 316 -656
rect 309 -661 648 -657
rect -436 -739 -418 -735
rect -436 -744 -432 -739
rect 312 -744 316 -661
rect 1069 -735 1073 -549
rect 1069 -739 1101 -735
rect 1069 -744 1073 -739
rect -436 -748 1073 -744
<< m5contact >>
rect 336 -64 341 -59
rect 360 -241 365 -236
rect 332 -410 337 -405
<< metal5 >>
rect 336 -237 340 -64
rect 336 -241 360 -237
rect 336 -405 340 -241
rect 337 -410 340 -405
<< labels >>
rlabel metal1 0 42 4 46 1 b0
rlabel metal1 0 50 4 54 1 a0
rlabel metal2 296 67 300 71 1 p0
rlabel metal2 296 -82 300 -78 1 p1
rlabel metal2 296 -232 300 -228 1 p2
rlabel metal2 296 -381 300 -377 1 p3
rlabel metal2 296 -531 300 -527 1 p4
rlabel metal1 277 -27 281 -23 1 g0
rlabel metal1 277 -176 281 -172 1 g1
rlabel metal1 276 -326 280 -322 1 g2
rlabel metal1 276 -475 280 -471 1 g3
rlabel metal1 276 -625 280 -621 1 g4
rlabel metal2 1053 -33 1057 -29 1 s1
rlabel metal2 1053 -142 1057 -138 1 s2
rlabel metal2 1053 -252 1057 -248 1 s3
rlabel metal2 1053 -363 1057 -359 1 s4
rlabel metal3 -10 -14 -7 66 3 vdd
rlabel metal1 596 -550 600 -546 1 c5
rlabel metal1 0 -99 4 -95 1 a1
rlabel metal1 0 -107 4 -103 1 b1
rlabel metal1 0 -249 4 -245 1 a2
rlabel metal1 0 -257 4 -253 1 b2
rlabel metal1 0 -398 4 -394 1 a3
rlabel metal1 0 -406 4 -402 1 b3
rlabel metal1 0 -548 4 -544 1 a4
rlabel metal1 0 -556 4 -552 1 b4
rlabel metal2 -405 75 -401 79 1 da0
rlabel metal2 -204 74 -200 78 1 db0
rlabel metal2 -404 -118 -400 -114 1 da1
rlabel metal2 -406 -306 -402 -302 1 da2
rlabel metal2 -405 -497 -401 -493 1 da3
rlabel metal2 -403 -687 -399 -683 1 da4
rlabel metal2 -202 -688 -198 -684 1 db4
rlabel metal2 -204 -498 -200 -494 1 db3
rlabel metal2 -205 -307 -201 -303 1 db2
rlabel metal2 -203 -119 -199 -115 1 db1
rlabel metal4 722 -748 792 -744 1 gnd
rlabel metal1 530 73 533 76 1 S0_out
rlabel metal1 1273 72 1277 76 1 S1_out
rlabel metal1 1274 -121 1278 -117 1 S2_out
rlabel metal1 1272 -309 1276 -305 1 S3_out
rlabel metal1 1273 -500 1277 -496 1 S4_out
rlabel metal1 1275 -690 1279 -686 1 Cout_ff
rlabel metal2 1295 -560 1314 -556 1 clk
<< end >>
